module t1 (output reg signed v);

always @* v = 1;

endmodule
