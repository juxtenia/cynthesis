module bitcount( input clk, input rst, input start, input [31:0] in, output reg finish, output reg signed [31:0] bitcount);
reg signed [31:0] output_output_34;
reg [31:0] output_in_34;
reg signed [31:0] output_i_34;
reg control_34_follow;
wire control_34_end;
reg control_34_start;
wire signed [31:0] input_i_34;
wire signed [31:0] input_output_34;
wire [31:0] input_in_34;
reg signed [31:0] output_i_33;
reg [31:0] output_in_33;
reg signed [31:0] output_output_33;
reg control_33_follow;
wire control_33_end;
reg control_33_start;
wire signed [31:0] input_i_33;
wire signed [31:0] input_output_33;
wire [31:0] input_in_33;
reg signed [31:0] output_i_30;
reg signed [31:0] output_output_30;
reg [31:0] output_in_30;
wire [31:0] operation_30_20;
reg control_30_follow;
wire control_30_end;
reg control_30_start;
wire signed [31:0] input_i_30;
wire signed [31:0] input_output_30;
wire [31:0] input_in_30;
wire signed [31:0] return_29;
reg control_29_follow;
wire control_29_end;
wire control_29_start;
wire signed [31:0] input_output_29;
reg signed [31:0] output_i_24;
reg signed [31:0] output_output_24;
reg [31:0] output_in_24;
wire signed [31:0] operation_24_11;
reg control_24_follow;
wire control_24_end;
reg control_24_start;
wire signed [31:0] input_i_24;
wire signed [31:0] input_output_24;
wire [31:0] input_in_24;
wire [31:0] output_in_20;
wire signed [31:0] output_output_20;
wire signed [31:0] output_i_20;
reg control_20_follow;
wire control_20_end;
wire control_20_start;
wire [31:0] input_in_20;
reg startfollow;

    assign input_i_34 = ((control_30_follow)?(output_i_30):((control_33_follow)?(output_i_33):(1'd0)));
    assign input_output_34 = ((control_30_follow)?(output_output_30):((control_33_follow)?(output_output_33):(1'd0)));
    assign input_in_34 = ((control_30_follow)?(output_in_30):((control_33_follow)?(output_in_33):(1'd0)));
    assign input_i_33 = (output_i_30);
    assign input_output_33 = (output_output_30);
    assign input_in_33 = (output_in_30);
    assign input_i_30 = (output_i_24);
    assign input_output_30 = (output_output_24);
    assign input_in_30 = (output_in_24);
    assign input_output_29 = (output_output_24);
    assign control_29_start = ((control_24_end)&&(!(operation_24_11)));
    assign input_i_24 = ((control_20_follow)?(output_i_20):((control_34_follow)?(output_i_34):(1'd0)));
    assign input_output_24 = ((control_20_follow)?(output_output_20):((control_34_follow)?(output_output_34):(1'd0)));
    assign input_in_24 = ((control_20_follow)?(output_in_20):((control_34_follow)?(output_in_34):(1'd0)));
    assign input_in_20 = (in);
    assign control_20_start = ((start)&&(!(startfollow)));
    assign control_34_end = (control_34_start);
    assign control_33_end = (control_33_start);
    assign operation_30_20 = ((input_in_30)&((32'd1)<<(input_i_30)));
    assign control_30_end = (control_30_start);
    assign return_29 = (input_output_29);
    assign control_29_end = (control_29_start);
    assign operation_24_11 = ((input_i_24)<(64'd32));
    assign control_24_end = (control_24_start);
    assign output_in_20 = (input_in_20);
    assign output_output_20 = (32'd0);
    assign output_i_20 = (32'd0);
    assign control_20_end = (control_20_start);
    
    always_ff @(posedge clk)
    if(rst)
         begin
            finish <= 1'd0;
            bitcount <= 32'd0;
            output_output_34 <= 32'd0;
            output_in_34 <= 32'd0;
            output_i_34 <= 32'd0;
            control_34_follow <= 1'd0;
            control_34_start <= 1'd0;
            output_i_33 <= 32'd0;
            output_in_33 <= 32'd0;
            output_output_33 <= 32'd0;
            control_33_follow <= 1'd0;
            control_33_start <= 1'd0;
            output_i_30 <= 32'd0;
            output_output_30 <= 32'd0;
            output_in_30 <= 32'd0;
            control_30_follow <= 1'd0;
            control_30_start <= 1'd0;
            control_29_follow <= 1'd0;
            output_i_24 <= 32'd0;
            output_output_24 <= 32'd0;
            output_in_24 <= 32'd0;
            control_24_follow <= 1'd0;
            control_24_start <= 1'd0;
            control_20_follow <= 1'd0;
            startfollow <= 1'd0;
        end
    else
        begin
            bitcount <= ((control_29_follow)?(return_29):(bitcount));
            finish <= ((!((start)&&(!(startfollow))))&&((finish)||(control_29_end)));
            control_34_start <= (((1'd0)||(control_33_end))||((control_30_end)&&(!(operation_30_20))));
            control_33_start <= ((control_30_end)&&(operation_30_20));
            control_30_start <= ((control_24_end)&&(operation_24_11));
            control_24_start <= (((1'd0)||(control_34_end))||(control_20_end));
            output_output_34 <= (input_output_34);
            output_in_34 <= (input_in_34);
            output_i_34 <= ((input_i_34)+(32'd1));
            control_34_follow <= (control_34_end);
            output_i_33 <= (input_i_33);
            output_in_33 <= (input_in_33);
            output_output_33 <= ((input_output_33)+(32'd1));
            control_33_follow <= (control_33_end);
            output_i_30 <= (input_i_30);
            output_output_30 <= (input_output_30);
            output_in_30 <= (input_in_30);
            control_30_follow <= (control_30_end);
            control_29_follow = (control_29_end);
            output_i_24 <= (input_i_24);
            output_output_24 <= (input_output_24);
            output_in_24 <= (input_in_24);
            control_24_follow <= (control_24_end);
            control_20_follow = (control_20_end);
            startfollow <= (start);
        end
endmodule // end of module bitcount
