module addkey( input clk, input rst, input start, input [127:0] in, input [127:0] key, output reg finish, output reg [127:0] addkey);
wire [127:0] return_186;
wire [7:0] operation_186_127;
reg signed [31:0] operation_186_126;
wire signed [31:0] operation_186_123;
wire [7:0] operation_186_7;
reg signed [31:0] operation_186_6;
wire [7:0] operation_186_23;
reg signed [31:0] operation_186_22;
wire [7:0] operation_186_39;
reg signed [31:0] operation_186_38;
wire [7:0] operation_186_55;
reg signed [31:0] operation_186_54;
wire [7:0] operation_186_71;
reg signed [31:0] operation_186_70;
wire [7:0] operation_186_87;
reg signed [31:0] operation_186_86;
wire [7:0] operation_186_103;
reg signed [31:0] operation_186_102;
wire [7:0] operation_186_119;
reg signed [31:0] operation_186_118;
wire signed [31:0] operation_186_117;
wire signed [31:0] operation_186_115;
wire signed [31:0] operation_186_101;
wire signed [31:0] operation_186_99;
wire signed [31:0] operation_186_85;
wire signed [31:0] operation_186_83;
wire signed [31:0] operation_186_69;
wire signed [31:0] operation_186_67;
wire signed [31:0] operation_186_53;
wire signed [31:0] operation_186_51;
wire signed [31:0] operation_186_37;
wire signed [31:0] operation_186_35;
wire signed [31:0] operation_186_21;
wire signed [31:0] operation_186_19;
wire signed [31:0] operation_186_5;
wire signed [31:0] operation_186_3;
wire [7:0] operation_186_15;
reg signed [31:0] operation_186_14;
wire signed [31:0] operation_186_11;
wire signed [31:0] operation_186_13;
wire [7:0] operation_186_31;
reg signed [31:0] operation_186_30;
wire signed [31:0] operation_186_27;
wire signed [31:0] operation_186_29;
wire [7:0] operation_186_47;
reg signed [31:0] operation_186_46;
wire signed [31:0] operation_186_43;
wire signed [31:0] operation_186_45;
wire [7:0] operation_186_63;
reg signed [31:0] operation_186_62;
wire signed [31:0] operation_186_59;
wire signed [31:0] operation_186_61;
wire [7:0] operation_186_79;
reg signed [31:0] operation_186_78;
wire signed [31:0] operation_186_75;
wire signed [31:0] operation_186_77;
wire [7:0] operation_186_95;
reg signed [31:0] operation_186_94;
wire signed [31:0] operation_186_91;
wire signed [31:0] operation_186_93;
wire [7:0] operation_186_111;
reg signed [31:0] operation_186_110;
wire signed [31:0] operation_186_107;
wire signed [31:0] operation_186_109;
wire signed [31:0] operation_186_125;
wire [127:0] operation_186_122;
wire [127:0] operation_186_124;
reg control_186_follow;
wire control_186_end;
wire control_186_0;
reg control_186_start;
reg [127:0] input_in_186_follow;
wire [127:0] input_in_186;
reg [127:0] input_key_186_follow;
wire [127:0] input_key_186;
reg startfollow;
initial begin
    
    
end
    assign input_in_186 = ((start)?(in):(input_in_186_follow));
    assign input_key_186 = ((start)?(key):(input_key_186_follow));
    assign return_186 = ({(operation_186_7[7:0]),(operation_186_15[7:0]),(operation_186_23[7:0]),(operation_186_31[7:0]),(operation_186_39[7:0]),(operation_186_47[7:0]),(operation_186_55[7:0]),(operation_186_63[7:0]),(operation_186_71[7:0]),(operation_186_79[7:0]),(operation_186_87[7:0]),(operation_186_95[7:0]),(operation_186_103[7:0]),(operation_186_111[7:0]),(operation_186_119[7:0]),(operation_186_127[7:0])});
    assign operation_186_127 = (operation_186_126);
    assign operation_186_123 = ({(operation_186_122[127:120])});
    assign operation_186_7 = (operation_186_6);
    assign operation_186_23 = (operation_186_22);
    assign operation_186_39 = (operation_186_38);
    assign operation_186_55 = (operation_186_54);
    assign operation_186_71 = (operation_186_70);
    assign operation_186_87 = (operation_186_86);
    assign operation_186_103 = (operation_186_102);
    assign operation_186_119 = (operation_186_118);
    assign operation_186_117 = ({(operation_186_124[119:112])});
    assign operation_186_115 = ({(operation_186_122[119:112])});
    assign operation_186_101 = ({(operation_186_124[103:96])});
    assign operation_186_99 = ({(operation_186_122[103:96])});
    assign operation_186_85 = ({(operation_186_124[87:80])});
    assign operation_186_83 = ({(operation_186_122[87:80])});
    assign operation_186_69 = ({(operation_186_124[71:64])});
    assign operation_186_67 = ({(operation_186_122[71:64])});
    assign operation_186_53 = ({(operation_186_124[55:48])});
    assign operation_186_51 = ({(operation_186_122[55:48])});
    assign operation_186_37 = ({(operation_186_124[39:32])});
    assign operation_186_35 = ({(operation_186_122[39:32])});
    assign operation_186_21 = ({(operation_186_124[23:16])});
    assign operation_186_19 = ({(operation_186_122[23:16])});
    assign operation_186_5 = ({(operation_186_124[7:0])});
    assign operation_186_3 = ({(operation_186_122[7:0])});
    assign operation_186_15 = (operation_186_14);
    assign operation_186_11 = ({(operation_186_122[15:8])});
    assign operation_186_13 = ({(operation_186_124[15:8])});
    assign operation_186_31 = (operation_186_30);
    assign operation_186_27 = ({(operation_186_122[31:24])});
    assign operation_186_29 = ({(operation_186_124[31:24])});
    assign operation_186_47 = (operation_186_46);
    assign operation_186_43 = ({(operation_186_122[47:40])});
    assign operation_186_45 = ({(operation_186_124[47:40])});
    assign operation_186_63 = (operation_186_62);
    assign operation_186_59 = ({(operation_186_122[63:56])});
    assign operation_186_61 = ({(operation_186_124[63:56])});
    assign operation_186_79 = (operation_186_78);
    assign operation_186_75 = ({(operation_186_122[79:72])});
    assign operation_186_77 = ({(operation_186_124[79:72])});
    assign operation_186_95 = (operation_186_94);
    assign operation_186_91 = ({(operation_186_122[95:88])});
    assign operation_186_93 = ({(operation_186_124[95:88])});
    assign operation_186_111 = (operation_186_110);
    assign operation_186_107 = ({(operation_186_122[111:104])});
    assign operation_186_109 = ({(operation_186_124[111:104])});
    assign operation_186_125 = ({(operation_186_124[127:120])});
    assign operation_186_122 = (input_in_186);
    assign operation_186_124 = (input_key_186);
    assign control_186_end = (control_186_start);
    assign control_186_0 = (control_186_start);
    
    always_ff @(posedge clk)
    if(rst)
         begin
            finish <= 1'd0;
            addkey <= 128'd0;
            operation_186_126 <= 32'd0;
            operation_186_6 <= 32'd0;
            operation_186_22 <= 32'd0;
            operation_186_38 <= 32'd0;
            operation_186_54 <= 32'd0;
            operation_186_70 <= 32'd0;
            operation_186_86 <= 32'd0;
            operation_186_102 <= 32'd0;
            operation_186_118 <= 32'd0;
            operation_186_14 <= 32'd0;
            operation_186_30 <= 32'd0;
            operation_186_46 <= 32'd0;
            operation_186_62 <= 32'd0;
            operation_186_78 <= 32'd0;
            operation_186_94 <= 32'd0;
            operation_186_110 <= 32'd0;
            control_186_follow <= 1'd0;
            control_186_start <= 1'd0;
            input_in_186_follow <= 128'd0;
            input_key_186_follow <= 128'd0;
            startfollow <= 1'd0;
        end
    else
        begin
            addkey <= ((control_186_follow)?(return_186):(addkey));
            finish <= ((!((start)&&(!(startfollow))))&&((finish)||(control_186_end)));
            control_186_start <= ((start)&&(!(startfollow)));
            operation_186_126 <= ((operation_186_123)^(operation_186_125));
            operation_186_6 <= ((operation_186_3)^(operation_186_5));
            operation_186_22 <= ((operation_186_19)^(operation_186_21));
            operation_186_38 <= ((operation_186_35)^(operation_186_37));
            operation_186_54 <= ((operation_186_51)^(operation_186_53));
            operation_186_70 <= ((operation_186_67)^(operation_186_69));
            operation_186_86 <= ((operation_186_83)^(operation_186_85));
            operation_186_102 <= ((operation_186_99)^(operation_186_101));
            operation_186_118 <= ((operation_186_115)^(operation_186_117));
            operation_186_14 <= ((operation_186_11)^(operation_186_13));
            operation_186_30 <= ((operation_186_27)^(operation_186_29));
            operation_186_46 <= ((operation_186_43)^(operation_186_45));
            operation_186_62 <= ((operation_186_59)^(operation_186_61));
            operation_186_78 <= ((operation_186_75)^(operation_186_77));
            operation_186_94 <= ((operation_186_91)^(operation_186_93));
            operation_186_110 <= ((operation_186_107)^(operation_186_109));
            control_186_follow <= (control_186_end);
            input_in_186_follow <= (input_in_186);
            input_key_186_follow <= (input_key_186);
            startfollow <= (start);
        end
endmodule // end of module addkey
