module AES128_encrypt( input clk, input rst, input start, input [127:0] in, input [127:0] key, output reg finish, output reg [127:0] AES128_encrypt);
wire [127:0] return_194;
wire [7:0] operation_194_1665;
reg signed [31:0] operation_194_1664;
wire signed [31:0] operation_194_1663;
wire [7:0] operation_194_1537;
reg signed [31:0] operation_194_1536;
wire [7:0] operation_194_1633;
wire [7:0] operation_194_1681;
reg signed [31:0] operation_194_1680;
wire signed [31:0] operation_194_1679;
reg signed [31:0] operation_194_1632;
wire signed [31:0] operation_194_1535;
wire [7:0] operation_194_1673;
reg signed [31:0] operation_194_1672;
wire [7:0] operation_194_1689;
reg signed [31:0] operation_194_1688;
wire signed [31:0] operation_194_1687;
wire signed [31:0] operation_194_1671;
wire [7:0] operation_194_1505;
reg signed [31:0] operation_194_1504;
wire [7:0] operation_194_1553;
reg signed [31:0] operation_194_1552;
wire [7:0] operation_194_1601;
wire [7:0] operation_194_1649;
reg signed [31:0] operation_194_1648;
reg signed [31:0] operation_194_1600;
wire signed [31:0] operation_194_1551;
wire signed [31:0] operation_194_1503;
wire [7:0] operation_194_1545;
reg signed [31:0] operation_194_1544;
wire [7:0] operation_194_1561;
reg signed [31:0] operation_194_1560;
wire [7:0] operation_194_1641;
wire [7:0] operation_194_1657;
reg signed [31:0] operation_194_1656;
reg signed [31:0] operation_194_1640;
wire signed [31:0] operation_194_1559;
wire signed [31:0] operation_194_1543;
wire [7:0] operation_194_1473;
reg signed [31:0] operation_194_1472;
wire [7:0] operation_194_1521;
reg signed [31:0] operation_194_1520;
wire [7:0] operation_194_1569;
wire [7:0] operation_194_1617;
reg signed [31:0] operation_194_1616;
reg signed [31:0] operation_194_1568;
wire signed [31:0] operation_194_1519;
wire signed [31:0] operation_194_1471;
wire [7:0] operation_194_1513;
reg signed [31:0] operation_194_1512;
wire [7:0] operation_194_1529;
reg signed [31:0] operation_194_1528;
wire [7:0] operation_194_1609;
wire [7:0] operation_194_1625;
reg signed [31:0] operation_194_1624;
reg signed [31:0] operation_194_1608;
wire signed [31:0] operation_194_1527;
wire signed [31:0] operation_194_1511;
wire [7:0] operation_194_1441;
reg signed [31:0] operation_194_1440;
wire [7:0] operation_194_1489;
reg signed [31:0] operation_194_1488;
wire [7:0] operation_194_1585;
reg signed [31:0] operation_194_1584;
wire signed [31:0] operation_194_1487;
wire signed [31:0] operation_194_1439;
wire [7:0] operation_194_1433;
reg signed [31:0] operation_194_1432;
wire [7:0] operation_194_1481;
reg signed [31:0] operation_194_1480;
wire [7:0] operation_194_1497;
reg signed [31:0] operation_194_1496;
wire [7:0] operation_194_1577;
wire [7:0] operation_194_1593;
reg signed [31:0] operation_194_1592;
reg signed [31:0] operation_194_1576;
wire signed [31:0] operation_194_1495;
wire signed [31:0] operation_194_1479;
wire signed [31:0] operation_194_1428;
wire [7:0] operation_194_1457;
reg signed [31:0] operation_194_1456;
wire signed [31:0] operation_194_1455;
wire [7:0] operation_194_1449;
reg signed [31:0] operation_194_1448;
wire [7:0] operation_194_1465;
reg signed [31:0] operation_194_1464;
wire signed [31:0] operation_194_1685;
wire signed [31:0] operation_194_1669;
wire signed [31:0] operation_194_1653;
wire signed [31:0] operation_194_1637;
wire signed [31:0] operation_194_1621;
wire signed [31:0] operation_194_1605;
wire signed [31:0] operation_194_1589;
wire signed [31:0] operation_194_1573;
wire signed [31:0] operation_194_1463;
wire signed [31:0] operation_194_1447;
wire signed [31:0] operation_194_1677;
wire signed [31:0] operation_194_1661;
wire signed [31:0] operation_194_1645;
wire signed [31:0] operation_194_1629;
wire signed [31:0] operation_194_1613;
wire signed [31:0] operation_194_1597;
wire signed [31:0] operation_194_1581;
wire signed [31:0] operation_194_1565;
reg [7:0] operation_194_1338_latch;
wire [7:0] operation_194_1338;
reg [7:0] operation_194_1328_latch;
wire [7:0] operation_194_1328;
reg [7:0] operation_194_1318_latch;
wire [7:0] operation_194_1318;
reg [7:0] operation_194_1308_latch;
wire [7:0] operation_194_1308;
reg [7:0] operation_194_1298_latch;
wire [7:0] operation_194_1298;
reg [7:0] operation_194_1288_latch;
wire [7:0] operation_194_1288;
reg [7:0] operation_194_1278_latch;
wire [7:0] operation_194_1278;
reg [7:0] operation_194_1268_latch;
wire [7:0] operation_194_1268;
reg [7:0] operation_194_1273_latch;
wire [7:0] operation_194_1273;
reg [7:0] operation_194_1283_latch;
wire [7:0] operation_194_1283;
reg [7:0] operation_194_1293_latch;
wire [7:0] operation_194_1293;
reg [7:0] operation_194_1303_latch;
wire [7:0] operation_194_1303;
reg [7:0] operation_194_1313_latch;
wire [7:0] operation_194_1313;
reg [7:0] operation_194_1323_latch;
wire [7:0] operation_194_1323;
reg [7:0] operation_194_1333_latch;
wire [7:0] operation_194_1333;
reg [7:0] operation_194_1343_latch;
wire [7:0] operation_194_1343;
reg [7:0] operation_194_1413_latch;
wire [7:0] operation_194_1413;
reg [7:0] operation_194_1423_latch;
wire [7:0] operation_194_1423;
reg [7:0] operation_194_1408_latch;
wire [7:0] operation_194_1408;
reg [7:0] operation_194_1418_latch;
wire [7:0] operation_194_1418;
wire [7:0] operation_194_5131;
reg signed [31:0] operation_194_5132;
wire signed [31:0] operation_194_5133;
wire [7:0] operation_194_5135;
reg signed [31:0] operation_194_5136;
wire [7:0] operation_194_5137;
reg signed [31:0] operation_194_5138;
wire [7:0] operation_194_5139;
reg signed [31:0] operation_194_5140;
wire [7:0] operation_194_5141;
reg signed [31:0] operation_194_5142;
wire [7:0] operation_194_5143;
reg signed [31:0] operation_194_5144;
wire [7:0] operation_194_5145;
reg signed [31:0] operation_194_5146;
wire [7:0] operation_194_5147;
reg signed [31:0] operation_194_5148;
wire [7:0] operation_194_5149;
reg signed [31:0] operation_194_5150;
wire signed [31:0] operation_194_5151;
wire signed [31:0] operation_194_5152;
wire signed [31:0] operation_194_5153;
wire signed [31:0] operation_194_5154;
wire signed [31:0] operation_194_5155;
wire signed [31:0] operation_194_5156;
wire signed [31:0] operation_194_5157;
wire signed [31:0] operation_194_5158;
wire signed [31:0] operation_194_5159;
wire signed [31:0] operation_194_5160;
wire [7:0] operation_194_5161;
reg signed [31:0] operation_194_5162;
wire [7:0] operation_194_5163;
reg signed [31:0] operation_194_5164;
wire [7:0] operation_194_5165;
reg signed [31:0] operation_194_5166;
wire [7:0] operation_194_5167;
reg signed [31:0] operation_194_5168;
wire [7:0] operation_194_5169;
reg signed [31:0] operation_194_5170;
wire [7:0] operation_194_5171;
reg signed [31:0] operation_194_5172;
wire [7:0] operation_194_5173;
reg signed [31:0] operation_194_5174;
wire [7:0] operation_194_5175;
reg signed [31:0] operation_194_5176;
wire [7:0] operation_194_5177;
reg signed [31:0] operation_194_5178;
wire [7:0] operation_194_5179;
reg signed [31:0] operation_194_5180;
wire [7:0] operation_194_5181;
reg signed [31:0] operation_194_5182;
wire [7:0] operation_194_5183;
reg signed [31:0] operation_194_5184;
wire [7:0] operation_194_5185;
reg signed [31:0] operation_194_5186;
wire [7:0] operation_194_5187;
reg signed [31:0] operation_194_5188;
wire [7:0] operation_194_5189;
reg signed [31:0] operation_194_5190;
wire [7:0] operation_194_5191;
reg signed [31:0] operation_194_5192;
wire signed [31:0] operation_194_5193;
wire signed [31:0] operation_194_5194;
wire signed [31:0] operation_194_5195;
wire signed [31:0] operation_194_5196;
wire signed [31:0] operation_194_5197;
wire signed [31:0] operation_194_5198;
wire signed [31:0] operation_194_5199;
wire signed [31:0] operation_194_5200;
wire signed [31:0] operation_194_5201;
wire signed [31:0] operation_194_5202;
wire signed [31:0] operation_194_5203;
wire signed [31:0] operation_194_5204;
wire signed [31:0] operation_194_5205;
wire signed [31:0] operation_194_5206;
wire signed [31:0] operation_194_5207;
wire signed [31:0] operation_194_5208;
wire signed [31:0] operation_194_5209;
wire signed [31:0] operation_194_5210;
wire [7:0] operation_194_5211;
reg signed [31:0] operation_194_5212;
wire [7:0] operation_194_5213;
reg signed [31:0] operation_194_5214;
wire [7:0] operation_194_5215;
reg signed [31:0] operation_194_5216;
wire [7:0] operation_194_5217;
reg signed [31:0] operation_194_5218;
wire [7:0] operation_194_5219;
reg signed [31:0] operation_194_5220;
wire [7:0] operation_194_5221;
reg signed [31:0] operation_194_5222;
wire [7:0] operation_194_5223;
reg signed [31:0] operation_194_5224;
wire [7:0] operation_194_5225;
reg signed [31:0] operation_194_5226;
wire [7:0] operation_194_5227;
reg signed [31:0] operation_194_5228;
wire [7:0] operation_194_5229;
reg signed [31:0] operation_194_5230;
wire signed [31:0] operation_194_5231;
wire signed [31:0] operation_194_5232;
wire signed [31:0] operation_194_5233;
wire signed [31:0] operation_194_5234;
wire signed [31:0] operation_194_5235;
wire signed [31:0] operation_194_5236;
wire signed [31:0] operation_194_5237;
wire signed [31:0] operation_194_5238;
wire signed [31:0] operation_194_5239;
wire signed [31:0] operation_194_5240;
wire [7:0] operation_194_5241;
reg signed [31:0] operation_194_5242;
wire [7:0] operation_194_5243;
reg signed [31:0] operation_194_5244;
wire [7:0] operation_194_5245;
reg signed [31:0] operation_194_5246;
wire [7:0] operation_194_5247;
reg signed [31:0] operation_194_5248;
wire [7:0] operation_194_5249;
reg signed [31:0] operation_194_5250;
wire [7:0] operation_194_5251;
reg signed [31:0] operation_194_5252;
wire [7:0] operation_194_5253;
reg signed [31:0] operation_194_5254;
wire [7:0] operation_194_5255;
reg signed [31:0] operation_194_5256;
wire [7:0] operation_194_5257;
reg signed [31:0] operation_194_5258;
wire [7:0] operation_194_5259;
reg signed [31:0] operation_194_5260;
wire signed [31:0] operation_194_5261;
wire signed [31:0] operation_194_5262;
wire signed [31:0] operation_194_5263;
wire signed [31:0] operation_194_5264;
wire signed [31:0] operation_194_5265;
wire signed [31:0] operation_194_5266;
wire signed [31:0] operation_194_5267;
wire signed [31:0] operation_194_5268;
wire signed [31:0] operation_194_5269;
wire signed [31:0] operation_194_5270;
wire [7:0] operation_194_5271;
reg signed [31:0] operation_194_5272;
wire [7:0] operation_194_5273;
reg signed [31:0] operation_194_5274;
wire [7:0] operation_194_5275;
reg signed [31:0] operation_194_5276;
wire [7:0] operation_194_5277;
reg signed [31:0] operation_194_5278;
wire [7:0] operation_194_5279;
reg signed [31:0] operation_194_5280;
wire [7:0] operation_194_5281;
reg signed [31:0] operation_194_5282;
wire [7:0] operation_194_5283;
reg signed [31:0] operation_194_5284;
wire [7:0] operation_194_5285;
reg signed [31:0] operation_194_5286;
wire [7:0] operation_194_5287;
reg signed [31:0] operation_194_5288;
wire [7:0] operation_194_5289;
reg signed [31:0] operation_194_5290;
wire signed [31:0] operation_194_5291;
wire signed [31:0] operation_194_5292;
wire signed [31:0] operation_194_5293;
wire signed [31:0] operation_194_5294;
wire signed [31:0] operation_194_5295;
wire signed [31:0] operation_194_5296;
wire signed [31:0] operation_194_5297;
wire signed [31:0] operation_194_5298;
wire signed [31:0] operation_194_5299;
wire signed [31:0] operation_194_5300;
wire [7:0] operation_194_5301;
reg signed [31:0] operation_194_5302;
reg signed [31:0] operation_194_5303;
wire [7:0] operation_194_5304;
reg signed [31:0] operation_194_5305;
reg signed [31:0] operation_194_5306;
wire [7:0] operation_194_5307;
reg signed [31:0] operation_194_5308;
reg signed [31:0] operation_194_5309;
wire [7:0] operation_194_5310;
reg signed [31:0] operation_194_5311;
reg signed [31:0] operation_194_5312;
wire [7:0] operation_194_5313;
reg signed [31:0] operation_194_5314;
reg signed [31:0] operation_194_5315;
wire [7:0] operation_194_5316;
reg signed [31:0] operation_194_5317;
reg signed [31:0] operation_194_5318;
wire [7:0] operation_194_5319;
reg signed [31:0] operation_194_5320;
reg signed [31:0] operation_194_5321;
wire [7:0] operation_194_5322;
reg signed [31:0] operation_194_5323;
reg signed [31:0] operation_194_5324;
wire [7:0] operation_194_5325;
reg signed [31:0] operation_194_5326;
wire [7:0] operation_194_5327;
reg signed [31:0] operation_194_5328;
wire signed [31:0] operation_194_5329;
wire signed [31:0] operation_194_5330;
reg signed [31:0] operation_194_5331;
reg signed [31:0] operation_194_5332;
reg signed [31:0] operation_194_5333;
wire signed [31:0] operation_194_5334;
reg signed [31:0] operation_194_5335;
reg signed [31:0] operation_194_5336;
reg signed [31:0] operation_194_5337;
wire signed [31:0] operation_194_5338;
reg signed [31:0] operation_194_5339;
reg signed [31:0] operation_194_5340;
reg signed [31:0] operation_194_5341;
wire signed [31:0] operation_194_5342;
reg signed [31:0] operation_194_5343;
reg signed [31:0] operation_194_5344;
reg signed [31:0] operation_194_5345;
wire signed [31:0] operation_194_5346;
reg signed [31:0] operation_194_5347;
reg signed [31:0] operation_194_5348;
reg signed [31:0] operation_194_5349;
wire signed [31:0] operation_194_5350;
reg signed [31:0] operation_194_5351;
reg signed [31:0] operation_194_5352;
reg signed [31:0] operation_194_5353;
wire signed [31:0] operation_194_5354;
reg signed [31:0] operation_194_5355;
reg signed [31:0] operation_194_5356;
reg signed [31:0] operation_194_5357;
wire signed [31:0] operation_194_5358;
reg signed [31:0] operation_194_5359;
reg signed [31:0] operation_194_5360;
reg signed [31:0] operation_194_5361;
wire signed [31:0] operation_194_5362;
wire [7:0] operation_194_5363;
reg signed [31:0] operation_194_5364;
reg signed [31:0] operation_194_5365;
wire [7:0] operation_194_5366;
reg signed [31:0] operation_194_5367;
reg signed [31:0] operation_194_5368;
wire [7:0] operation_194_5369;
reg signed [31:0] operation_194_5370;
reg signed [31:0] operation_194_5371;
wire [7:0] operation_194_5372;
reg signed [31:0] operation_194_5373;
reg signed [31:0] operation_194_5374;
wire [7:0] operation_194_5375;
reg signed [31:0] operation_194_5376;
reg signed [31:0] operation_194_5377;
wire [7:0] operation_194_5378;
reg signed [31:0] operation_194_5379;
reg signed [31:0] operation_194_5380;
wire [7:0] operation_194_5381;
reg signed [31:0] operation_194_5382;
reg signed [31:0] operation_194_5383;
wire [7:0] operation_194_5384;
reg signed [31:0] operation_194_5385;
reg signed [31:0] operation_194_5386;
wire [7:0] operation_194_5387;
reg signed [31:0] operation_194_5388;
wire [7:0] operation_194_5389;
reg signed [31:0] operation_194_5390;
wire signed [31:0] operation_194_5391;
wire signed [31:0] operation_194_5392;
wire signed [31:0] operation_194_5393;
wire signed [31:0] operation_194_5394;
reg signed [31:0] operation_194_5395;
reg signed [31:0] operation_194_5396;
reg signed [31:0] operation_194_5397;
wire signed [31:0] operation_194_5398;
reg signed [31:0] operation_194_5399;
reg signed [31:0] operation_194_5400;
reg signed [31:0] operation_194_5401;
wire signed [31:0] operation_194_5402;
reg signed [31:0] operation_194_5403;
reg signed [31:0] operation_194_5404;
reg signed [31:0] operation_194_5405;
wire signed [31:0] operation_194_5406;
reg signed [31:0] operation_194_5407;
reg signed [31:0] operation_194_5408;
reg signed [31:0] operation_194_5409;
wire signed [31:0] operation_194_5410;
reg signed [31:0] operation_194_5411;
reg signed [31:0] operation_194_5412;
reg signed [31:0] operation_194_5413;
wire signed [31:0] operation_194_5414;
reg signed [31:0] operation_194_5415;
reg signed [31:0] operation_194_5416;
reg signed [31:0] operation_194_5417;
wire signed [31:0] operation_194_5418;
reg signed [31:0] operation_194_5419;
reg signed [31:0] operation_194_5420;
reg signed [31:0] operation_194_5421;
wire signed [31:0] operation_194_5422;
reg signed [31:0] operation_194_5423;
reg signed [31:0] operation_194_5424;
reg signed [31:0] operation_194_5425;
wire signed [31:0] operation_194_5426;
wire [7:0] operation_194_5427;
wire [7:0] operation_194_5428;
reg signed [31:0] operation_194_5429;
wire [7:0] operation_194_5430;
wire [7:0] operation_194_5431;
reg signed [31:0] operation_194_5432;
wire [7:0] operation_194_5433;
wire [7:0] operation_194_5434;
reg signed [31:0] operation_194_5435;
wire [7:0] operation_194_5436;
wire [7:0] operation_194_5437;
reg signed [31:0] operation_194_5438;
wire [7:0] operation_194_5439;
reg signed [31:0] operation_194_5440;
wire [7:0] operation_194_5441;
reg signed [31:0] operation_194_5442;
wire [7:0] operation_194_5443;
reg signed [31:0] operation_194_5444;
wire [7:0] operation_194_5445;
reg signed [31:0] operation_194_5446;
wire [7:0] operation_194_5447;
reg signed [31:0] operation_194_5448;
wire signed [31:0] operation_194_5449;
wire signed [31:0] operation_194_5450;
wire signed [31:0] operation_194_5451;
wire signed [31:0] operation_194_5452;
wire signed [31:0] operation_194_5453;
reg signed [31:0] operation_194_5454;
reg signed [31:0] operation_194_5455;
reg signed [31:0] operation_194_5456;
reg signed [31:0] operation_194_5457;
wire [7:0] operation_194_5458;
reg signed [31:0] operation_194_5459;
wire [7:0] operation_194_5460;
reg signed [31:0] operation_194_5461;
wire [7:0] operation_194_5462;
reg signed [31:0] operation_194_5463;
wire [7:0] operation_194_5464;
reg signed [31:0] operation_194_5465;
wire [7:0] operation_194_5466;
reg signed [31:0] operation_194_5467;
wire [7:0] operation_194_5468;
reg signed [31:0] operation_194_5469;
wire [7:0] operation_194_5470;
reg signed [31:0] operation_194_5471;
wire [7:0] operation_194_5472;
reg signed [31:0] operation_194_5473;
wire [7:0] operation_194_5474;
reg signed [31:0] operation_194_5475;
wire [7:0] operation_194_5476;
reg signed [31:0] operation_194_5477;
wire [7:0] operation_194_5478;
reg signed [31:0] operation_194_5479;
wire signed [31:0] operation_194_5486;
reg signed [31:0] operation_194_5489;
reg signed [31:0] operation_194_5490;
reg signed [31:0] operation_194_5491;
reg signed [31:0] operation_194_5492;
wire signed [31:0] operation_194_5493;
wire signed [31:0] operation_194_5494;
wire signed [31:0] operation_194_5495;
wire signed [31:0] operation_194_5496;
wire signed [31:0] operation_194_5497;
wire signed [31:0] operation_194_5498;
wire signed [31:0] operation_194_5499;
wire signed [31:0] operation_194_5500;
wire [7:0] operation_194_5503;
reg signed [31:0] operation_194_5504;
wire [7:0] operation_194_5505;
reg signed [31:0] operation_194_5506;
wire signed [31:0] operation_194_5517;
wire signed [31:0] operation_194_5519;
reg [7:0] operation_194_5521_latch;
wire [7:0] operation_194_5521;
reg [7:0] operation_194_5522_latch;
wire [7:0] operation_194_5522;
wire signed [31:0] operation_194_5523;
wire signed [31:0] operation_194_5524;
wire signed [31:0] operation_194_5525;
wire signed [31:0] operation_194_5526;
wire signed [31:0] operation_194_5527;
wire signed [31:0] operation_194_5528;
wire signed [31:0] operation_194_5529;
wire signed [31:0] operation_194_5530;
reg [7:0] operation_194_5531_latch;
wire [7:0] operation_194_5531;
reg [7:0] operation_194_5532_latch;
wire [7:0] operation_194_5532;
reg [7:0] operation_194_5533_latch;
wire [7:0] operation_194_5533;
reg [7:0] operation_194_5534_latch;
wire [7:0] operation_194_5534;
reg [7:0] operation_194_5535_latch;
wire [7:0] operation_194_5535;
reg [7:0] operation_194_5536_latch;
wire [7:0] operation_194_5536;
reg [7:0] operation_194_5537_latch;
wire [7:0] operation_194_5537;
reg [7:0] operation_194_5538_latch;
wire [7:0] operation_194_5538;
reg [7:0] operation_194_5539_latch;
wire [7:0] operation_194_5539;
reg [7:0] operation_194_5540_latch;
wire [7:0] operation_194_5540;
reg [7:0] operation_194_5541_latch;
wire [7:0] operation_194_5541;
reg [7:0] operation_194_5542_latch;
wire [7:0] operation_194_5542;
reg [7:0] operation_194_5543_latch;
wire [7:0] operation_194_5543;
reg [7:0] operation_194_5544_latch;
wire [7:0] operation_194_5544;
reg [7:0] operation_194_5545_latch;
wire [7:0] operation_194_5545;
reg [7:0] operation_194_5546_latch;
wire [7:0] operation_194_5546;
reg [7:0] operation_194_5547_latch;
wire [7:0] operation_194_5547;
reg [7:0] operation_194_5548_latch;
wire [7:0] operation_194_5548;
wire [7:0] operation_194_4702;
reg signed [31:0] operation_194_4703;
wire signed [31:0] operation_194_4704;
wire [7:0] operation_194_4706;
reg signed [31:0] operation_194_4707;
wire [7:0] operation_194_4708;
reg signed [31:0] operation_194_4709;
wire [7:0] operation_194_4710;
reg signed [31:0] operation_194_4711;
wire [7:0] operation_194_4712;
reg signed [31:0] operation_194_4713;
wire [7:0] operation_194_4714;
reg signed [31:0] operation_194_4715;
wire [7:0] operation_194_4716;
reg signed [31:0] operation_194_4717;
wire [7:0] operation_194_4718;
reg signed [31:0] operation_194_4719;
wire [7:0] operation_194_4720;
reg signed [31:0] operation_194_4721;
wire signed [31:0] operation_194_4722;
wire signed [31:0] operation_194_4723;
wire signed [31:0] operation_194_4724;
wire signed [31:0] operation_194_4725;
wire signed [31:0] operation_194_4726;
wire signed [31:0] operation_194_4727;
wire signed [31:0] operation_194_4728;
wire signed [31:0] operation_194_4729;
wire signed [31:0] operation_194_4730;
wire signed [31:0] operation_194_4731;
wire [7:0] operation_194_4732;
reg signed [31:0] operation_194_4733;
wire [7:0] operation_194_4734;
reg signed [31:0] operation_194_4735;
wire [7:0] operation_194_4736;
reg signed [31:0] operation_194_4737;
wire [7:0] operation_194_4738;
reg signed [31:0] operation_194_4739;
wire [7:0] operation_194_4740;
reg signed [31:0] operation_194_4741;
wire [7:0] operation_194_4742;
reg signed [31:0] operation_194_4743;
wire [7:0] operation_194_4744;
reg signed [31:0] operation_194_4745;
wire [7:0] operation_194_4746;
reg signed [31:0] operation_194_4747;
wire [7:0] operation_194_4748;
reg signed [31:0] operation_194_4749;
wire [7:0] operation_194_4750;
reg signed [31:0] operation_194_4751;
wire [7:0] operation_194_4752;
reg signed [31:0] operation_194_4753;
wire [7:0] operation_194_4754;
reg signed [31:0] operation_194_4755;
wire [7:0] operation_194_4756;
reg signed [31:0] operation_194_4757;
wire [7:0] operation_194_4758;
reg signed [31:0] operation_194_4759;
wire [7:0] operation_194_4760;
reg signed [31:0] operation_194_4761;
wire [7:0] operation_194_4762;
reg signed [31:0] operation_194_4763;
wire signed [31:0] operation_194_4764;
wire signed [31:0] operation_194_4765;
wire signed [31:0] operation_194_4766;
wire signed [31:0] operation_194_4767;
wire signed [31:0] operation_194_4768;
wire signed [31:0] operation_194_4769;
wire signed [31:0] operation_194_4770;
wire signed [31:0] operation_194_4771;
wire signed [31:0] operation_194_4772;
wire signed [31:0] operation_194_4773;
wire signed [31:0] operation_194_4774;
wire signed [31:0] operation_194_4775;
wire signed [31:0] operation_194_4776;
wire signed [31:0] operation_194_4777;
wire signed [31:0] operation_194_4778;
wire signed [31:0] operation_194_4779;
wire signed [31:0] operation_194_4780;
wire signed [31:0] operation_194_4781;
wire [7:0] operation_194_4782;
reg signed [31:0] operation_194_4783;
wire [7:0] operation_194_4784;
reg signed [31:0] operation_194_4785;
wire [7:0] operation_194_4786;
reg signed [31:0] operation_194_4787;
wire [7:0] operation_194_4788;
reg signed [31:0] operation_194_4789;
wire [7:0] operation_194_4790;
reg signed [31:0] operation_194_4791;
wire [7:0] operation_194_4792;
reg signed [31:0] operation_194_4793;
wire [7:0] operation_194_4794;
reg signed [31:0] operation_194_4795;
wire [7:0] operation_194_4796;
reg signed [31:0] operation_194_4797;
wire [7:0] operation_194_4798;
reg signed [31:0] operation_194_4799;
wire [7:0] operation_194_4800;
reg signed [31:0] operation_194_4801;
wire signed [31:0] operation_194_4802;
wire signed [31:0] operation_194_4803;
wire signed [31:0] operation_194_4804;
wire signed [31:0] operation_194_4805;
wire signed [31:0] operation_194_4806;
wire signed [31:0] operation_194_4807;
wire signed [31:0] operation_194_4808;
wire signed [31:0] operation_194_4809;
wire signed [31:0] operation_194_4810;
wire signed [31:0] operation_194_4811;
wire [7:0] operation_194_4812;
reg signed [31:0] operation_194_4813;
wire [7:0] operation_194_4814;
reg signed [31:0] operation_194_4815;
wire [7:0] operation_194_4816;
reg signed [31:0] operation_194_4817;
wire [7:0] operation_194_4818;
reg signed [31:0] operation_194_4819;
wire [7:0] operation_194_4820;
reg signed [31:0] operation_194_4821;
wire [7:0] operation_194_4822;
reg signed [31:0] operation_194_4823;
wire [7:0] operation_194_4824;
reg signed [31:0] operation_194_4825;
wire [7:0] operation_194_4826;
reg signed [31:0] operation_194_4827;
wire [7:0] operation_194_4828;
reg signed [31:0] operation_194_4829;
wire [7:0] operation_194_4830;
reg signed [31:0] operation_194_4831;
wire signed [31:0] operation_194_4832;
wire signed [31:0] operation_194_4833;
wire signed [31:0] operation_194_4834;
wire signed [31:0] operation_194_4835;
wire signed [31:0] operation_194_4836;
wire signed [31:0] operation_194_4837;
wire signed [31:0] operation_194_4838;
wire signed [31:0] operation_194_4839;
wire signed [31:0] operation_194_4840;
wire signed [31:0] operation_194_4841;
wire [7:0] operation_194_4842;
reg signed [31:0] operation_194_4843;
wire [7:0] operation_194_4844;
reg signed [31:0] operation_194_4845;
wire [7:0] operation_194_4846;
reg signed [31:0] operation_194_4847;
wire [7:0] operation_194_4848;
reg signed [31:0] operation_194_4849;
wire [7:0] operation_194_4850;
reg signed [31:0] operation_194_4851;
wire [7:0] operation_194_4852;
reg signed [31:0] operation_194_4853;
wire [7:0] operation_194_4854;
reg signed [31:0] operation_194_4855;
wire [7:0] operation_194_4856;
reg signed [31:0] operation_194_4857;
wire [7:0] operation_194_4858;
reg signed [31:0] operation_194_4859;
wire [7:0] operation_194_4860;
reg signed [31:0] operation_194_4861;
wire signed [31:0] operation_194_4862;
wire signed [31:0] operation_194_4863;
wire signed [31:0] operation_194_4864;
wire signed [31:0] operation_194_4865;
wire signed [31:0] operation_194_4866;
wire signed [31:0] operation_194_4867;
wire signed [31:0] operation_194_4868;
wire signed [31:0] operation_194_4869;
wire signed [31:0] operation_194_4870;
wire signed [31:0] operation_194_4871;
wire [7:0] operation_194_4872;
reg signed [31:0] operation_194_4873;
reg signed [31:0] operation_194_4874;
wire [7:0] operation_194_4875;
reg signed [31:0] operation_194_4876;
reg signed [31:0] operation_194_4877;
wire [7:0] operation_194_4878;
reg signed [31:0] operation_194_4879;
reg signed [31:0] operation_194_4880;
wire [7:0] operation_194_4881;
reg signed [31:0] operation_194_4882;
reg signed [31:0] operation_194_4883;
wire [7:0] operation_194_4884;
reg signed [31:0] operation_194_4885;
reg signed [31:0] operation_194_4886;
wire [7:0] operation_194_4887;
reg signed [31:0] operation_194_4888;
reg signed [31:0] operation_194_4889;
wire [7:0] operation_194_4890;
reg signed [31:0] operation_194_4891;
reg signed [31:0] operation_194_4892;
wire [7:0] operation_194_4893;
reg signed [31:0] operation_194_4894;
reg signed [31:0] operation_194_4895;
wire [7:0] operation_194_4896;
reg signed [31:0] operation_194_4897;
wire [7:0] operation_194_4898;
reg signed [31:0] operation_194_4899;
wire signed [31:0] operation_194_4900;
wire signed [31:0] operation_194_4901;
reg signed [31:0] operation_194_4902;
reg signed [31:0] operation_194_4903;
reg signed [31:0] operation_194_4904;
wire signed [31:0] operation_194_4905;
reg signed [31:0] operation_194_4906;
reg signed [31:0] operation_194_4907;
reg signed [31:0] operation_194_4908;
wire signed [31:0] operation_194_4909;
reg signed [31:0] operation_194_4910;
reg signed [31:0] operation_194_4911;
reg signed [31:0] operation_194_4912;
wire signed [31:0] operation_194_4913;
reg signed [31:0] operation_194_4914;
reg signed [31:0] operation_194_4915;
reg signed [31:0] operation_194_4916;
wire signed [31:0] operation_194_4917;
reg signed [31:0] operation_194_4918;
reg signed [31:0] operation_194_4919;
reg signed [31:0] operation_194_4920;
wire signed [31:0] operation_194_4921;
reg signed [31:0] operation_194_4922;
reg signed [31:0] operation_194_4923;
reg signed [31:0] operation_194_4924;
wire signed [31:0] operation_194_4925;
reg signed [31:0] operation_194_4926;
reg signed [31:0] operation_194_4927;
reg signed [31:0] operation_194_4928;
wire signed [31:0] operation_194_4929;
reg signed [31:0] operation_194_4930;
reg signed [31:0] operation_194_4931;
reg signed [31:0] operation_194_4932;
wire signed [31:0] operation_194_4933;
wire [7:0] operation_194_4934;
reg signed [31:0] operation_194_4935;
reg signed [31:0] operation_194_4936;
wire [7:0] operation_194_4937;
reg signed [31:0] operation_194_4938;
reg signed [31:0] operation_194_4939;
wire [7:0] operation_194_4940;
reg signed [31:0] operation_194_4941;
reg signed [31:0] operation_194_4942;
wire [7:0] operation_194_4943;
reg signed [31:0] operation_194_4944;
reg signed [31:0] operation_194_4945;
wire [7:0] operation_194_4946;
reg signed [31:0] operation_194_4947;
reg signed [31:0] operation_194_4948;
wire [7:0] operation_194_4949;
reg signed [31:0] operation_194_4950;
reg signed [31:0] operation_194_4951;
wire [7:0] operation_194_4952;
reg signed [31:0] operation_194_4953;
reg signed [31:0] operation_194_4954;
wire [7:0] operation_194_4955;
reg signed [31:0] operation_194_4956;
reg signed [31:0] operation_194_4957;
wire [7:0] operation_194_4958;
reg signed [31:0] operation_194_4959;
wire [7:0] operation_194_4960;
reg signed [31:0] operation_194_4961;
wire signed [31:0] operation_194_4962;
wire signed [31:0] operation_194_4963;
wire signed [31:0] operation_194_4964;
wire signed [31:0] operation_194_4965;
reg signed [31:0] operation_194_4966;
reg signed [31:0] operation_194_4967;
reg signed [31:0] operation_194_4968;
wire signed [31:0] operation_194_4969;
reg signed [31:0] operation_194_4970;
reg signed [31:0] operation_194_4971;
reg signed [31:0] operation_194_4972;
wire signed [31:0] operation_194_4973;
reg signed [31:0] operation_194_4974;
reg signed [31:0] operation_194_4975;
reg signed [31:0] operation_194_4976;
wire signed [31:0] operation_194_4977;
reg signed [31:0] operation_194_4978;
reg signed [31:0] operation_194_4979;
reg signed [31:0] operation_194_4980;
wire signed [31:0] operation_194_4981;
reg signed [31:0] operation_194_4982;
reg signed [31:0] operation_194_4983;
reg signed [31:0] operation_194_4984;
wire signed [31:0] operation_194_4985;
reg signed [31:0] operation_194_4986;
reg signed [31:0] operation_194_4987;
reg signed [31:0] operation_194_4988;
wire signed [31:0] operation_194_4989;
reg signed [31:0] operation_194_4990;
reg signed [31:0] operation_194_4991;
reg signed [31:0] operation_194_4992;
wire signed [31:0] operation_194_4993;
reg signed [31:0] operation_194_4994;
reg signed [31:0] operation_194_4995;
reg signed [31:0] operation_194_4996;
wire signed [31:0] operation_194_4997;
wire [7:0] operation_194_4998;
wire [7:0] operation_194_4999;
reg signed [31:0] operation_194_5000;
wire [7:0] operation_194_5001;
wire [7:0] operation_194_5002;
reg signed [31:0] operation_194_5003;
wire [7:0] operation_194_5004;
wire [7:0] operation_194_5005;
reg signed [31:0] operation_194_5006;
wire [7:0] operation_194_5007;
wire [7:0] operation_194_5008;
reg signed [31:0] operation_194_5009;
wire [7:0] operation_194_5010;
reg signed [31:0] operation_194_5011;
wire [7:0] operation_194_5012;
reg signed [31:0] operation_194_5013;
wire [7:0] operation_194_5014;
reg signed [31:0] operation_194_5015;
wire [7:0] operation_194_5016;
reg signed [31:0] operation_194_5017;
wire [7:0] operation_194_5018;
reg signed [31:0] operation_194_5019;
wire signed [31:0] operation_194_5020;
wire signed [31:0] operation_194_5021;
wire signed [31:0] operation_194_5022;
wire signed [31:0] operation_194_5023;
wire signed [31:0] operation_194_5024;
reg signed [31:0] operation_194_5025;
reg signed [31:0] operation_194_5026;
reg signed [31:0] operation_194_5027;
reg signed [31:0] operation_194_5028;
wire [7:0] operation_194_5029;
reg signed [31:0] operation_194_5030;
wire [7:0] operation_194_5031;
reg signed [31:0] operation_194_5032;
wire [7:0] operation_194_5033;
reg signed [31:0] operation_194_5034;
wire [7:0] operation_194_5035;
reg signed [31:0] operation_194_5036;
wire [7:0] operation_194_5037;
reg signed [31:0] operation_194_5038;
wire [7:0] operation_194_5039;
reg signed [31:0] operation_194_5040;
wire [7:0] operation_194_5041;
reg signed [31:0] operation_194_5042;
wire [7:0] operation_194_5043;
reg signed [31:0] operation_194_5044;
wire [7:0] operation_194_5045;
reg signed [31:0] operation_194_5046;
wire [7:0] operation_194_5047;
reg signed [31:0] operation_194_5048;
wire [7:0] operation_194_5049;
reg signed [31:0] operation_194_5050;
wire signed [31:0] operation_194_5057;
reg signed [31:0] operation_194_5060;
reg signed [31:0] operation_194_5061;
reg signed [31:0] operation_194_5062;
reg signed [31:0] operation_194_5063;
wire signed [31:0] operation_194_5064;
wire signed [31:0] operation_194_5065;
wire signed [31:0] operation_194_5066;
wire signed [31:0] operation_194_5067;
wire signed [31:0] operation_194_5068;
wire signed [31:0] operation_194_5069;
wire signed [31:0] operation_194_5070;
wire signed [31:0] operation_194_5071;
wire [7:0] operation_194_5074;
reg signed [31:0] operation_194_5075;
wire [7:0] operation_194_5076;
reg signed [31:0] operation_194_5077;
wire signed [31:0] operation_194_5088;
wire signed [31:0] operation_194_5090;
reg [7:0] operation_194_5092_latch;
wire [7:0] operation_194_5092;
reg [7:0] operation_194_5093_latch;
wire [7:0] operation_194_5093;
wire signed [31:0] operation_194_5094;
wire signed [31:0] operation_194_5095;
wire signed [31:0] operation_194_5096;
wire signed [31:0] operation_194_5097;
wire signed [31:0] operation_194_5098;
wire signed [31:0] operation_194_5099;
wire signed [31:0] operation_194_5100;
wire signed [31:0] operation_194_5101;
reg [7:0] operation_194_5102_latch;
wire [7:0] operation_194_5102;
reg [7:0] operation_194_5103_latch;
wire [7:0] operation_194_5103;
reg [7:0] operation_194_5104_latch;
wire [7:0] operation_194_5104;
reg [7:0] operation_194_5105_latch;
wire [7:0] operation_194_5105;
reg [7:0] operation_194_5106_latch;
wire [7:0] operation_194_5106;
reg [7:0] operation_194_5107_latch;
wire [7:0] operation_194_5107;
reg [7:0] operation_194_5108_latch;
wire [7:0] operation_194_5108;
reg [7:0] operation_194_5109_latch;
wire [7:0] operation_194_5109;
reg [7:0] operation_194_5110_latch;
wire [7:0] operation_194_5110;
reg [7:0] operation_194_5111_latch;
wire [7:0] operation_194_5111;
reg [7:0] operation_194_5112_latch;
wire [7:0] operation_194_5112;
reg [7:0] operation_194_5113_latch;
wire [7:0] operation_194_5113;
reg [7:0] operation_194_5114_latch;
wire [7:0] operation_194_5114;
reg [7:0] operation_194_5115_latch;
wire [7:0] operation_194_5115;
reg [7:0] operation_194_5116_latch;
wire [7:0] operation_194_5116;
reg [7:0] operation_194_5117_latch;
wire [7:0] operation_194_5117;
reg [7:0] operation_194_5118_latch;
wire [7:0] operation_194_5118;
reg [7:0] operation_194_5119_latch;
wire [7:0] operation_194_5119;
wire [7:0] operation_194_4273;
reg signed [31:0] operation_194_4274;
wire signed [31:0] operation_194_4275;
wire [7:0] operation_194_4277;
reg signed [31:0] operation_194_4278;
wire [7:0] operation_194_4279;
reg signed [31:0] operation_194_4280;
wire [7:0] operation_194_4281;
reg signed [31:0] operation_194_4282;
wire [7:0] operation_194_4283;
reg signed [31:0] operation_194_4284;
wire [7:0] operation_194_4285;
reg signed [31:0] operation_194_4286;
wire [7:0] operation_194_4287;
reg signed [31:0] operation_194_4288;
wire [7:0] operation_194_4289;
reg signed [31:0] operation_194_4290;
wire [7:0] operation_194_4291;
reg signed [31:0] operation_194_4292;
wire signed [31:0] operation_194_4293;
wire signed [31:0] operation_194_4294;
wire signed [31:0] operation_194_4295;
wire signed [31:0] operation_194_4296;
wire signed [31:0] operation_194_4297;
wire signed [31:0] operation_194_4298;
wire signed [31:0] operation_194_4299;
wire signed [31:0] operation_194_4300;
wire signed [31:0] operation_194_4301;
wire signed [31:0] operation_194_4302;
wire [7:0] operation_194_4303;
reg signed [31:0] operation_194_4304;
wire [7:0] operation_194_4305;
reg signed [31:0] operation_194_4306;
wire [7:0] operation_194_4307;
reg signed [31:0] operation_194_4308;
wire [7:0] operation_194_4309;
reg signed [31:0] operation_194_4310;
wire [7:0] operation_194_4311;
reg signed [31:0] operation_194_4312;
wire [7:0] operation_194_4313;
reg signed [31:0] operation_194_4314;
wire [7:0] operation_194_4315;
reg signed [31:0] operation_194_4316;
wire [7:0] operation_194_4317;
reg signed [31:0] operation_194_4318;
wire [7:0] operation_194_4319;
reg signed [31:0] operation_194_4320;
wire [7:0] operation_194_4321;
reg signed [31:0] operation_194_4322;
wire [7:0] operation_194_4323;
reg signed [31:0] operation_194_4324;
wire [7:0] operation_194_4325;
reg signed [31:0] operation_194_4326;
wire [7:0] operation_194_4327;
reg signed [31:0] operation_194_4328;
wire [7:0] operation_194_4329;
reg signed [31:0] operation_194_4330;
wire [7:0] operation_194_4331;
reg signed [31:0] operation_194_4332;
wire [7:0] operation_194_4333;
reg signed [31:0] operation_194_4334;
wire signed [31:0] operation_194_4335;
wire signed [31:0] operation_194_4336;
wire signed [31:0] operation_194_4337;
wire signed [31:0] operation_194_4338;
wire signed [31:0] operation_194_4339;
wire signed [31:0] operation_194_4340;
wire signed [31:0] operation_194_4341;
wire signed [31:0] operation_194_4342;
wire signed [31:0] operation_194_4343;
wire signed [31:0] operation_194_4344;
wire signed [31:0] operation_194_4345;
wire signed [31:0] operation_194_4346;
wire signed [31:0] operation_194_4347;
wire signed [31:0] operation_194_4348;
wire signed [31:0] operation_194_4349;
wire signed [31:0] operation_194_4350;
wire signed [31:0] operation_194_4351;
wire signed [31:0] operation_194_4352;
wire [7:0] operation_194_4353;
reg signed [31:0] operation_194_4354;
wire [7:0] operation_194_4355;
reg signed [31:0] operation_194_4356;
wire [7:0] operation_194_4357;
reg signed [31:0] operation_194_4358;
wire [7:0] operation_194_4359;
reg signed [31:0] operation_194_4360;
wire [7:0] operation_194_4361;
reg signed [31:0] operation_194_4362;
wire [7:0] operation_194_4363;
reg signed [31:0] operation_194_4364;
wire [7:0] operation_194_4365;
reg signed [31:0] operation_194_4366;
wire [7:0] operation_194_4367;
reg signed [31:0] operation_194_4368;
wire [7:0] operation_194_4369;
reg signed [31:0] operation_194_4370;
wire [7:0] operation_194_4371;
reg signed [31:0] operation_194_4372;
wire signed [31:0] operation_194_4373;
wire signed [31:0] operation_194_4374;
wire signed [31:0] operation_194_4375;
wire signed [31:0] operation_194_4376;
wire signed [31:0] operation_194_4377;
wire signed [31:0] operation_194_4378;
wire signed [31:0] operation_194_4379;
wire signed [31:0] operation_194_4380;
wire signed [31:0] operation_194_4381;
wire signed [31:0] operation_194_4382;
wire [7:0] operation_194_4383;
reg signed [31:0] operation_194_4384;
wire [7:0] operation_194_4385;
reg signed [31:0] operation_194_4386;
wire [7:0] operation_194_4387;
reg signed [31:0] operation_194_4388;
wire [7:0] operation_194_4389;
reg signed [31:0] operation_194_4390;
wire [7:0] operation_194_4391;
reg signed [31:0] operation_194_4392;
wire [7:0] operation_194_4393;
reg signed [31:0] operation_194_4394;
wire [7:0] operation_194_4395;
reg signed [31:0] operation_194_4396;
wire [7:0] operation_194_4397;
reg signed [31:0] operation_194_4398;
wire [7:0] operation_194_4399;
reg signed [31:0] operation_194_4400;
wire [7:0] operation_194_4401;
reg signed [31:0] operation_194_4402;
wire signed [31:0] operation_194_4403;
wire signed [31:0] operation_194_4404;
wire signed [31:0] operation_194_4405;
wire signed [31:0] operation_194_4406;
wire signed [31:0] operation_194_4407;
wire signed [31:0] operation_194_4408;
wire signed [31:0] operation_194_4409;
wire signed [31:0] operation_194_4410;
wire signed [31:0] operation_194_4411;
wire signed [31:0] operation_194_4412;
wire [7:0] operation_194_4413;
reg signed [31:0] operation_194_4414;
wire [7:0] operation_194_4415;
reg signed [31:0] operation_194_4416;
wire [7:0] operation_194_4417;
reg signed [31:0] operation_194_4418;
wire [7:0] operation_194_4419;
reg signed [31:0] operation_194_4420;
wire [7:0] operation_194_4421;
reg signed [31:0] operation_194_4422;
wire [7:0] operation_194_4423;
reg signed [31:0] operation_194_4424;
wire [7:0] operation_194_4425;
reg signed [31:0] operation_194_4426;
wire [7:0] operation_194_4427;
reg signed [31:0] operation_194_4428;
wire [7:0] operation_194_4429;
reg signed [31:0] operation_194_4430;
wire [7:0] operation_194_4431;
reg signed [31:0] operation_194_4432;
wire signed [31:0] operation_194_4433;
wire signed [31:0] operation_194_4434;
wire signed [31:0] operation_194_4435;
wire signed [31:0] operation_194_4436;
wire signed [31:0] operation_194_4437;
wire signed [31:0] operation_194_4438;
wire signed [31:0] operation_194_4439;
wire signed [31:0] operation_194_4440;
wire signed [31:0] operation_194_4441;
wire signed [31:0] operation_194_4442;
wire [7:0] operation_194_4443;
reg signed [31:0] operation_194_4444;
reg signed [31:0] operation_194_4445;
wire [7:0] operation_194_4446;
reg signed [31:0] operation_194_4447;
reg signed [31:0] operation_194_4448;
wire [7:0] operation_194_4449;
reg signed [31:0] operation_194_4450;
reg signed [31:0] operation_194_4451;
wire [7:0] operation_194_4452;
reg signed [31:0] operation_194_4453;
reg signed [31:0] operation_194_4454;
wire [7:0] operation_194_4455;
reg signed [31:0] operation_194_4456;
reg signed [31:0] operation_194_4457;
wire [7:0] operation_194_4458;
reg signed [31:0] operation_194_4459;
reg signed [31:0] operation_194_4460;
wire [7:0] operation_194_4461;
reg signed [31:0] operation_194_4462;
reg signed [31:0] operation_194_4463;
wire [7:0] operation_194_4464;
reg signed [31:0] operation_194_4465;
reg signed [31:0] operation_194_4466;
wire [7:0] operation_194_4467;
reg signed [31:0] operation_194_4468;
wire [7:0] operation_194_4469;
reg signed [31:0] operation_194_4470;
wire signed [31:0] operation_194_4471;
wire signed [31:0] operation_194_4472;
reg signed [31:0] operation_194_4473;
reg signed [31:0] operation_194_4474;
reg signed [31:0] operation_194_4475;
wire signed [31:0] operation_194_4476;
reg signed [31:0] operation_194_4477;
reg signed [31:0] operation_194_4478;
reg signed [31:0] operation_194_4479;
wire signed [31:0] operation_194_4480;
reg signed [31:0] operation_194_4481;
reg signed [31:0] operation_194_4482;
reg signed [31:0] operation_194_4483;
wire signed [31:0] operation_194_4484;
reg signed [31:0] operation_194_4485;
reg signed [31:0] operation_194_4486;
reg signed [31:0] operation_194_4487;
wire signed [31:0] operation_194_4488;
reg signed [31:0] operation_194_4489;
reg signed [31:0] operation_194_4490;
reg signed [31:0] operation_194_4491;
wire signed [31:0] operation_194_4492;
reg signed [31:0] operation_194_4493;
reg signed [31:0] operation_194_4494;
reg signed [31:0] operation_194_4495;
wire signed [31:0] operation_194_4496;
reg signed [31:0] operation_194_4497;
reg signed [31:0] operation_194_4498;
reg signed [31:0] operation_194_4499;
wire signed [31:0] operation_194_4500;
reg signed [31:0] operation_194_4501;
reg signed [31:0] operation_194_4502;
reg signed [31:0] operation_194_4503;
wire signed [31:0] operation_194_4504;
wire [7:0] operation_194_4505;
reg signed [31:0] operation_194_4506;
reg signed [31:0] operation_194_4507;
wire [7:0] operation_194_4508;
reg signed [31:0] operation_194_4509;
reg signed [31:0] operation_194_4510;
wire [7:0] operation_194_4511;
reg signed [31:0] operation_194_4512;
reg signed [31:0] operation_194_4513;
wire [7:0] operation_194_4514;
reg signed [31:0] operation_194_4515;
reg signed [31:0] operation_194_4516;
wire [7:0] operation_194_4517;
reg signed [31:0] operation_194_4518;
reg signed [31:0] operation_194_4519;
wire [7:0] operation_194_4520;
reg signed [31:0] operation_194_4521;
reg signed [31:0] operation_194_4522;
wire [7:0] operation_194_4523;
reg signed [31:0] operation_194_4524;
reg signed [31:0] operation_194_4525;
wire [7:0] operation_194_4526;
reg signed [31:0] operation_194_4527;
reg signed [31:0] operation_194_4528;
wire [7:0] operation_194_4529;
reg signed [31:0] operation_194_4530;
wire [7:0] operation_194_4531;
reg signed [31:0] operation_194_4532;
wire signed [31:0] operation_194_4533;
wire signed [31:0] operation_194_4534;
wire signed [31:0] operation_194_4535;
wire signed [31:0] operation_194_4536;
reg signed [31:0] operation_194_4537;
reg signed [31:0] operation_194_4538;
reg signed [31:0] operation_194_4539;
wire signed [31:0] operation_194_4540;
reg signed [31:0] operation_194_4541;
reg signed [31:0] operation_194_4542;
reg signed [31:0] operation_194_4543;
wire signed [31:0] operation_194_4544;
reg signed [31:0] operation_194_4545;
reg signed [31:0] operation_194_4546;
reg signed [31:0] operation_194_4547;
wire signed [31:0] operation_194_4548;
reg signed [31:0] operation_194_4549;
reg signed [31:0] operation_194_4550;
reg signed [31:0] operation_194_4551;
wire signed [31:0] operation_194_4552;
reg signed [31:0] operation_194_4553;
reg signed [31:0] operation_194_4554;
reg signed [31:0] operation_194_4555;
wire signed [31:0] operation_194_4556;
reg signed [31:0] operation_194_4557;
reg signed [31:0] operation_194_4558;
reg signed [31:0] operation_194_4559;
wire signed [31:0] operation_194_4560;
reg signed [31:0] operation_194_4561;
reg signed [31:0] operation_194_4562;
reg signed [31:0] operation_194_4563;
wire signed [31:0] operation_194_4564;
reg signed [31:0] operation_194_4565;
reg signed [31:0] operation_194_4566;
reg signed [31:0] operation_194_4567;
wire signed [31:0] operation_194_4568;
wire [7:0] operation_194_4569;
wire [7:0] operation_194_4570;
reg signed [31:0] operation_194_4571;
wire [7:0] operation_194_4572;
wire [7:0] operation_194_4573;
reg signed [31:0] operation_194_4574;
wire [7:0] operation_194_4575;
wire [7:0] operation_194_4576;
reg signed [31:0] operation_194_4577;
wire [7:0] operation_194_4578;
wire [7:0] operation_194_4579;
reg signed [31:0] operation_194_4580;
wire [7:0] operation_194_4581;
reg signed [31:0] operation_194_4582;
wire [7:0] operation_194_4583;
reg signed [31:0] operation_194_4584;
wire [7:0] operation_194_4585;
reg signed [31:0] operation_194_4586;
wire [7:0] operation_194_4587;
reg signed [31:0] operation_194_4588;
wire [7:0] operation_194_4589;
reg signed [31:0] operation_194_4590;
wire signed [31:0] operation_194_4591;
wire signed [31:0] operation_194_4592;
wire signed [31:0] operation_194_4593;
wire signed [31:0] operation_194_4594;
wire signed [31:0] operation_194_4595;
reg signed [31:0] operation_194_4596;
reg signed [31:0] operation_194_4597;
reg signed [31:0] operation_194_4598;
reg signed [31:0] operation_194_4599;
wire [7:0] operation_194_4600;
reg signed [31:0] operation_194_4601;
wire [7:0] operation_194_4602;
reg signed [31:0] operation_194_4603;
wire [7:0] operation_194_4604;
reg signed [31:0] operation_194_4605;
wire [7:0] operation_194_4606;
reg signed [31:0] operation_194_4607;
wire [7:0] operation_194_4608;
reg signed [31:0] operation_194_4609;
wire [7:0] operation_194_4610;
reg signed [31:0] operation_194_4611;
wire [7:0] operation_194_4612;
reg signed [31:0] operation_194_4613;
wire [7:0] operation_194_4614;
reg signed [31:0] operation_194_4615;
wire [7:0] operation_194_4616;
reg signed [31:0] operation_194_4617;
wire [7:0] operation_194_4618;
reg signed [31:0] operation_194_4619;
wire [7:0] operation_194_4620;
reg signed [31:0] operation_194_4621;
wire signed [31:0] operation_194_4628;
reg signed [31:0] operation_194_4631;
reg signed [31:0] operation_194_4632;
reg signed [31:0] operation_194_4633;
reg signed [31:0] operation_194_4634;
wire signed [31:0] operation_194_4635;
wire signed [31:0] operation_194_4636;
wire signed [31:0] operation_194_4637;
wire signed [31:0] operation_194_4638;
wire signed [31:0] operation_194_4639;
wire signed [31:0] operation_194_4640;
wire signed [31:0] operation_194_4641;
wire signed [31:0] operation_194_4642;
wire [7:0] operation_194_4645;
reg signed [31:0] operation_194_4646;
wire [7:0] operation_194_4647;
reg signed [31:0] operation_194_4648;
wire signed [31:0] operation_194_4659;
wire signed [31:0] operation_194_4661;
reg [7:0] operation_194_4663_latch;
wire [7:0] operation_194_4663;
reg [7:0] operation_194_4664_latch;
wire [7:0] operation_194_4664;
wire signed [31:0] operation_194_4665;
wire signed [31:0] operation_194_4666;
wire signed [31:0] operation_194_4667;
wire signed [31:0] operation_194_4668;
wire signed [31:0] operation_194_4669;
wire signed [31:0] operation_194_4670;
wire signed [31:0] operation_194_4671;
wire signed [31:0] operation_194_4672;
reg [7:0] operation_194_4673_latch;
wire [7:0] operation_194_4673;
reg [7:0] operation_194_4674_latch;
wire [7:0] operation_194_4674;
reg [7:0] operation_194_4675_latch;
wire [7:0] operation_194_4675;
reg [7:0] operation_194_4676_latch;
wire [7:0] operation_194_4676;
reg [7:0] operation_194_4677_latch;
wire [7:0] operation_194_4677;
reg [7:0] operation_194_4678_latch;
wire [7:0] operation_194_4678;
reg [7:0] operation_194_4679_latch;
wire [7:0] operation_194_4679;
reg [7:0] operation_194_4680_latch;
wire [7:0] operation_194_4680;
reg [7:0] operation_194_4681_latch;
wire [7:0] operation_194_4681;
reg [7:0] operation_194_4682_latch;
wire [7:0] operation_194_4682;
reg [7:0] operation_194_4683_latch;
wire [7:0] operation_194_4683;
reg [7:0] operation_194_4684_latch;
wire [7:0] operation_194_4684;
reg [7:0] operation_194_4685_latch;
wire [7:0] operation_194_4685;
reg [7:0] operation_194_4686_latch;
wire [7:0] operation_194_4686;
reg [7:0] operation_194_4687_latch;
wire [7:0] operation_194_4687;
reg [7:0] operation_194_4688_latch;
wire [7:0] operation_194_4688;
reg [7:0] operation_194_4689_latch;
wire [7:0] operation_194_4689;
reg [7:0] operation_194_4690_latch;
wire [7:0] operation_194_4690;
wire [7:0] operation_194_3844;
reg signed [31:0] operation_194_3845;
wire signed [31:0] operation_194_3846;
wire [7:0] operation_194_3848;
reg signed [31:0] operation_194_3849;
wire [7:0] operation_194_3850;
reg signed [31:0] operation_194_3851;
wire [7:0] operation_194_3852;
reg signed [31:0] operation_194_3853;
wire [7:0] operation_194_3854;
reg signed [31:0] operation_194_3855;
wire [7:0] operation_194_3856;
reg signed [31:0] operation_194_3857;
wire [7:0] operation_194_3858;
reg signed [31:0] operation_194_3859;
wire [7:0] operation_194_3860;
reg signed [31:0] operation_194_3861;
wire [7:0] operation_194_3862;
reg signed [31:0] operation_194_3863;
wire signed [31:0] operation_194_3864;
wire signed [31:0] operation_194_3865;
wire signed [31:0] operation_194_3866;
wire signed [31:0] operation_194_3867;
wire signed [31:0] operation_194_3868;
wire signed [31:0] operation_194_3869;
wire signed [31:0] operation_194_3870;
wire signed [31:0] operation_194_3871;
wire signed [31:0] operation_194_3872;
wire signed [31:0] operation_194_3873;
wire [7:0] operation_194_3874;
reg signed [31:0] operation_194_3875;
wire [7:0] operation_194_3876;
reg signed [31:0] operation_194_3877;
wire [7:0] operation_194_3878;
reg signed [31:0] operation_194_3879;
wire [7:0] operation_194_3880;
reg signed [31:0] operation_194_3881;
wire [7:0] operation_194_3882;
reg signed [31:0] operation_194_3883;
wire [7:0] operation_194_3884;
reg signed [31:0] operation_194_3885;
wire [7:0] operation_194_3886;
reg signed [31:0] operation_194_3887;
wire [7:0] operation_194_3888;
reg signed [31:0] operation_194_3889;
wire [7:0] operation_194_3890;
reg signed [31:0] operation_194_3891;
wire [7:0] operation_194_3892;
reg signed [31:0] operation_194_3893;
wire [7:0] operation_194_3894;
reg signed [31:0] operation_194_3895;
wire [7:0] operation_194_3896;
reg signed [31:0] operation_194_3897;
wire [7:0] operation_194_3898;
reg signed [31:0] operation_194_3899;
wire [7:0] operation_194_3900;
reg signed [31:0] operation_194_3901;
wire [7:0] operation_194_3902;
reg signed [31:0] operation_194_3903;
wire [7:0] operation_194_3904;
reg signed [31:0] operation_194_3905;
wire signed [31:0] operation_194_3906;
wire signed [31:0] operation_194_3907;
wire signed [31:0] operation_194_3908;
wire signed [31:0] operation_194_3909;
wire signed [31:0] operation_194_3910;
wire signed [31:0] operation_194_3911;
wire signed [31:0] operation_194_3912;
wire signed [31:0] operation_194_3913;
wire signed [31:0] operation_194_3914;
wire signed [31:0] operation_194_3915;
wire signed [31:0] operation_194_3916;
wire signed [31:0] operation_194_3917;
wire signed [31:0] operation_194_3918;
wire signed [31:0] operation_194_3919;
wire signed [31:0] operation_194_3920;
wire signed [31:0] operation_194_3921;
wire signed [31:0] operation_194_3922;
wire signed [31:0] operation_194_3923;
wire [7:0] operation_194_3924;
reg signed [31:0] operation_194_3925;
wire [7:0] operation_194_3926;
reg signed [31:0] operation_194_3927;
wire [7:0] operation_194_3928;
reg signed [31:0] operation_194_3929;
wire [7:0] operation_194_3930;
reg signed [31:0] operation_194_3931;
wire [7:0] operation_194_3932;
reg signed [31:0] operation_194_3933;
wire [7:0] operation_194_3934;
reg signed [31:0] operation_194_3935;
wire [7:0] operation_194_3936;
reg signed [31:0] operation_194_3937;
wire [7:0] operation_194_3938;
reg signed [31:0] operation_194_3939;
wire [7:0] operation_194_3940;
reg signed [31:0] operation_194_3941;
wire [7:0] operation_194_3942;
reg signed [31:0] operation_194_3943;
wire signed [31:0] operation_194_3944;
wire signed [31:0] operation_194_3945;
wire signed [31:0] operation_194_3946;
wire signed [31:0] operation_194_3947;
wire signed [31:0] operation_194_3948;
wire signed [31:0] operation_194_3949;
wire signed [31:0] operation_194_3950;
wire signed [31:0] operation_194_3951;
wire signed [31:0] operation_194_3952;
wire signed [31:0] operation_194_3953;
wire [7:0] operation_194_3954;
reg signed [31:0] operation_194_3955;
wire [7:0] operation_194_3956;
reg signed [31:0] operation_194_3957;
wire [7:0] operation_194_3958;
reg signed [31:0] operation_194_3959;
wire [7:0] operation_194_3960;
reg signed [31:0] operation_194_3961;
wire [7:0] operation_194_3962;
reg signed [31:0] operation_194_3963;
wire [7:0] operation_194_3964;
reg signed [31:0] operation_194_3965;
wire [7:0] operation_194_3966;
reg signed [31:0] operation_194_3967;
wire [7:0] operation_194_3968;
reg signed [31:0] operation_194_3969;
wire [7:0] operation_194_3970;
reg signed [31:0] operation_194_3971;
wire [7:0] operation_194_3972;
reg signed [31:0] operation_194_3973;
wire signed [31:0] operation_194_3974;
wire signed [31:0] operation_194_3975;
wire signed [31:0] operation_194_3976;
wire signed [31:0] operation_194_3977;
wire signed [31:0] operation_194_3978;
wire signed [31:0] operation_194_3979;
wire signed [31:0] operation_194_3980;
wire signed [31:0] operation_194_3981;
wire signed [31:0] operation_194_3982;
wire signed [31:0] operation_194_3983;
wire [7:0] operation_194_3984;
reg signed [31:0] operation_194_3985;
wire [7:0] operation_194_3986;
reg signed [31:0] operation_194_3987;
wire [7:0] operation_194_3988;
reg signed [31:0] operation_194_3989;
wire [7:0] operation_194_3990;
reg signed [31:0] operation_194_3991;
wire [7:0] operation_194_3992;
reg signed [31:0] operation_194_3993;
wire [7:0] operation_194_3994;
reg signed [31:0] operation_194_3995;
wire [7:0] operation_194_3996;
reg signed [31:0] operation_194_3997;
wire [7:0] operation_194_3998;
reg signed [31:0] operation_194_3999;
wire [7:0] operation_194_4000;
reg signed [31:0] operation_194_4001;
wire [7:0] operation_194_4002;
reg signed [31:0] operation_194_4003;
wire signed [31:0] operation_194_4004;
wire signed [31:0] operation_194_4005;
wire signed [31:0] operation_194_4006;
wire signed [31:0] operation_194_4007;
wire signed [31:0] operation_194_4008;
wire signed [31:0] operation_194_4009;
wire signed [31:0] operation_194_4010;
wire signed [31:0] operation_194_4011;
wire signed [31:0] operation_194_4012;
wire signed [31:0] operation_194_4013;
wire [7:0] operation_194_4014;
reg signed [31:0] operation_194_4015;
reg signed [31:0] operation_194_4016;
wire [7:0] operation_194_4017;
reg signed [31:0] operation_194_4018;
reg signed [31:0] operation_194_4019;
wire [7:0] operation_194_4020;
reg signed [31:0] operation_194_4021;
reg signed [31:0] operation_194_4022;
wire [7:0] operation_194_4023;
reg signed [31:0] operation_194_4024;
reg signed [31:0] operation_194_4025;
wire [7:0] operation_194_4026;
reg signed [31:0] operation_194_4027;
reg signed [31:0] operation_194_4028;
wire [7:0] operation_194_4029;
reg signed [31:0] operation_194_4030;
reg signed [31:0] operation_194_4031;
wire [7:0] operation_194_4032;
reg signed [31:0] operation_194_4033;
reg signed [31:0] operation_194_4034;
wire [7:0] operation_194_4035;
reg signed [31:0] operation_194_4036;
reg signed [31:0] operation_194_4037;
wire [7:0] operation_194_4038;
reg signed [31:0] operation_194_4039;
wire [7:0] operation_194_4040;
reg signed [31:0] operation_194_4041;
wire signed [31:0] operation_194_4042;
wire signed [31:0] operation_194_4043;
reg signed [31:0] operation_194_4044;
reg signed [31:0] operation_194_4045;
reg signed [31:0] operation_194_4046;
wire signed [31:0] operation_194_4047;
reg signed [31:0] operation_194_4048;
reg signed [31:0] operation_194_4049;
reg signed [31:0] operation_194_4050;
wire signed [31:0] operation_194_4051;
reg signed [31:0] operation_194_4052;
reg signed [31:0] operation_194_4053;
reg signed [31:0] operation_194_4054;
wire signed [31:0] operation_194_4055;
reg signed [31:0] operation_194_4056;
reg signed [31:0] operation_194_4057;
reg signed [31:0] operation_194_4058;
wire signed [31:0] operation_194_4059;
reg signed [31:0] operation_194_4060;
reg signed [31:0] operation_194_4061;
reg signed [31:0] operation_194_4062;
wire signed [31:0] operation_194_4063;
reg signed [31:0] operation_194_4064;
reg signed [31:0] operation_194_4065;
reg signed [31:0] operation_194_4066;
wire signed [31:0] operation_194_4067;
reg signed [31:0] operation_194_4068;
reg signed [31:0] operation_194_4069;
reg signed [31:0] operation_194_4070;
wire signed [31:0] operation_194_4071;
reg signed [31:0] operation_194_4072;
reg signed [31:0] operation_194_4073;
reg signed [31:0] operation_194_4074;
wire signed [31:0] operation_194_4075;
wire [7:0] operation_194_4076;
reg signed [31:0] operation_194_4077;
reg signed [31:0] operation_194_4078;
wire [7:0] operation_194_4079;
reg signed [31:0] operation_194_4080;
reg signed [31:0] operation_194_4081;
wire [7:0] operation_194_4082;
reg signed [31:0] operation_194_4083;
reg signed [31:0] operation_194_4084;
wire [7:0] operation_194_4085;
reg signed [31:0] operation_194_4086;
reg signed [31:0] operation_194_4087;
wire [7:0] operation_194_4088;
reg signed [31:0] operation_194_4089;
reg signed [31:0] operation_194_4090;
wire [7:0] operation_194_4091;
reg signed [31:0] operation_194_4092;
reg signed [31:0] operation_194_4093;
wire [7:0] operation_194_4094;
reg signed [31:0] operation_194_4095;
reg signed [31:0] operation_194_4096;
wire [7:0] operation_194_4097;
reg signed [31:0] operation_194_4098;
reg signed [31:0] operation_194_4099;
wire [7:0] operation_194_4100;
reg signed [31:0] operation_194_4101;
wire [7:0] operation_194_4102;
reg signed [31:0] operation_194_4103;
wire signed [31:0] operation_194_4104;
wire signed [31:0] operation_194_4105;
wire signed [31:0] operation_194_4106;
wire signed [31:0] operation_194_4107;
reg signed [31:0] operation_194_4108;
reg signed [31:0] operation_194_4109;
reg signed [31:0] operation_194_4110;
wire signed [31:0] operation_194_4111;
reg signed [31:0] operation_194_4112;
reg signed [31:0] operation_194_4113;
reg signed [31:0] operation_194_4114;
wire signed [31:0] operation_194_4115;
reg signed [31:0] operation_194_4116;
reg signed [31:0] operation_194_4117;
reg signed [31:0] operation_194_4118;
wire signed [31:0] operation_194_4119;
reg signed [31:0] operation_194_4120;
reg signed [31:0] operation_194_4121;
reg signed [31:0] operation_194_4122;
wire signed [31:0] operation_194_4123;
reg signed [31:0] operation_194_4124;
reg signed [31:0] operation_194_4125;
reg signed [31:0] operation_194_4126;
wire signed [31:0] operation_194_4127;
reg signed [31:0] operation_194_4128;
reg signed [31:0] operation_194_4129;
reg signed [31:0] operation_194_4130;
wire signed [31:0] operation_194_4131;
reg signed [31:0] operation_194_4132;
reg signed [31:0] operation_194_4133;
reg signed [31:0] operation_194_4134;
wire signed [31:0] operation_194_4135;
reg signed [31:0] operation_194_4136;
reg signed [31:0] operation_194_4137;
reg signed [31:0] operation_194_4138;
wire signed [31:0] operation_194_4139;
wire [7:0] operation_194_4140;
wire [7:0] operation_194_4141;
reg signed [31:0] operation_194_4142;
wire [7:0] operation_194_4143;
wire [7:0] operation_194_4144;
reg signed [31:0] operation_194_4145;
wire [7:0] operation_194_4146;
wire [7:0] operation_194_4147;
reg signed [31:0] operation_194_4148;
wire [7:0] operation_194_4149;
wire [7:0] operation_194_4150;
reg signed [31:0] operation_194_4151;
wire [7:0] operation_194_4152;
reg signed [31:0] operation_194_4153;
wire [7:0] operation_194_4154;
reg signed [31:0] operation_194_4155;
wire [7:0] operation_194_4156;
reg signed [31:0] operation_194_4157;
wire [7:0] operation_194_4158;
reg signed [31:0] operation_194_4159;
wire [7:0] operation_194_4160;
reg signed [31:0] operation_194_4161;
wire signed [31:0] operation_194_4162;
wire signed [31:0] operation_194_4163;
wire signed [31:0] operation_194_4164;
wire signed [31:0] operation_194_4165;
wire signed [31:0] operation_194_4166;
reg signed [31:0] operation_194_4167;
reg signed [31:0] operation_194_4168;
reg signed [31:0] operation_194_4169;
reg signed [31:0] operation_194_4170;
wire [7:0] operation_194_4171;
reg signed [31:0] operation_194_4172;
wire [7:0] operation_194_4173;
reg signed [31:0] operation_194_4174;
wire [7:0] operation_194_4175;
reg signed [31:0] operation_194_4176;
wire [7:0] operation_194_4177;
reg signed [31:0] operation_194_4178;
wire [7:0] operation_194_4179;
reg signed [31:0] operation_194_4180;
wire [7:0] operation_194_4181;
reg signed [31:0] operation_194_4182;
wire [7:0] operation_194_4183;
reg signed [31:0] operation_194_4184;
wire [7:0] operation_194_4185;
reg signed [31:0] operation_194_4186;
wire [7:0] operation_194_4187;
reg signed [31:0] operation_194_4188;
wire [7:0] operation_194_4189;
reg signed [31:0] operation_194_4190;
wire [7:0] operation_194_4191;
reg signed [31:0] operation_194_4192;
wire signed [31:0] operation_194_4199;
reg signed [31:0] operation_194_4202;
reg signed [31:0] operation_194_4203;
reg signed [31:0] operation_194_4204;
reg signed [31:0] operation_194_4205;
wire signed [31:0] operation_194_4206;
wire signed [31:0] operation_194_4207;
wire signed [31:0] operation_194_4208;
wire signed [31:0] operation_194_4209;
wire signed [31:0] operation_194_4210;
wire signed [31:0] operation_194_4211;
wire signed [31:0] operation_194_4212;
wire signed [31:0] operation_194_4213;
wire [7:0] operation_194_4216;
reg signed [31:0] operation_194_4217;
wire [7:0] operation_194_4218;
reg signed [31:0] operation_194_4219;
wire signed [31:0] operation_194_4230;
wire signed [31:0] operation_194_4232;
reg [7:0] operation_194_4234_latch;
wire [7:0] operation_194_4234;
reg [7:0] operation_194_4235_latch;
wire [7:0] operation_194_4235;
wire signed [31:0] operation_194_4236;
wire signed [31:0] operation_194_4237;
wire signed [31:0] operation_194_4238;
wire signed [31:0] operation_194_4239;
wire signed [31:0] operation_194_4240;
wire signed [31:0] operation_194_4241;
wire signed [31:0] operation_194_4242;
wire signed [31:0] operation_194_4243;
reg [7:0] operation_194_4244_latch;
wire [7:0] operation_194_4244;
reg [7:0] operation_194_4245_latch;
wire [7:0] operation_194_4245;
reg [7:0] operation_194_4246_latch;
wire [7:0] operation_194_4246;
reg [7:0] operation_194_4247_latch;
wire [7:0] operation_194_4247;
reg [7:0] operation_194_4248_latch;
wire [7:0] operation_194_4248;
reg [7:0] operation_194_4249_latch;
wire [7:0] operation_194_4249;
reg [7:0] operation_194_4250_latch;
wire [7:0] operation_194_4250;
reg [7:0] operation_194_4251_latch;
wire [7:0] operation_194_4251;
reg [7:0] operation_194_4252_latch;
wire [7:0] operation_194_4252;
reg [7:0] operation_194_4253_latch;
wire [7:0] operation_194_4253;
reg [7:0] operation_194_4254_latch;
wire [7:0] operation_194_4254;
reg [7:0] operation_194_4255_latch;
wire [7:0] operation_194_4255;
reg [7:0] operation_194_4256_latch;
wire [7:0] operation_194_4256;
reg [7:0] operation_194_4257_latch;
wire [7:0] operation_194_4257;
reg [7:0] operation_194_4258_latch;
wire [7:0] operation_194_4258;
reg [7:0] operation_194_4259_latch;
wire [7:0] operation_194_4259;
reg [7:0] operation_194_4260_latch;
wire [7:0] operation_194_4260;
reg [7:0] operation_194_4261_latch;
wire [7:0] operation_194_4261;
wire [7:0] operation_194_3415;
reg signed [31:0] operation_194_3416;
wire signed [31:0] operation_194_3417;
wire [7:0] operation_194_3419;
reg signed [31:0] operation_194_3420;
wire [7:0] operation_194_3421;
reg signed [31:0] operation_194_3422;
wire [7:0] operation_194_3423;
reg signed [31:0] operation_194_3424;
wire [7:0] operation_194_3425;
reg signed [31:0] operation_194_3426;
wire [7:0] operation_194_3427;
reg signed [31:0] operation_194_3428;
wire [7:0] operation_194_3429;
reg signed [31:0] operation_194_3430;
wire [7:0] operation_194_3431;
reg signed [31:0] operation_194_3432;
wire [7:0] operation_194_3433;
reg signed [31:0] operation_194_3434;
wire signed [31:0] operation_194_3435;
wire signed [31:0] operation_194_3436;
wire signed [31:0] operation_194_3437;
wire signed [31:0] operation_194_3438;
wire signed [31:0] operation_194_3439;
wire signed [31:0] operation_194_3440;
wire signed [31:0] operation_194_3441;
wire signed [31:0] operation_194_3442;
wire signed [31:0] operation_194_3443;
wire signed [31:0] operation_194_3444;
wire [7:0] operation_194_3445;
reg signed [31:0] operation_194_3446;
wire [7:0] operation_194_3447;
reg signed [31:0] operation_194_3448;
wire [7:0] operation_194_3449;
reg signed [31:0] operation_194_3450;
wire [7:0] operation_194_3451;
reg signed [31:0] operation_194_3452;
wire [7:0] operation_194_3453;
reg signed [31:0] operation_194_3454;
wire [7:0] operation_194_3455;
reg signed [31:0] operation_194_3456;
wire [7:0] operation_194_3457;
reg signed [31:0] operation_194_3458;
wire [7:0] operation_194_3459;
reg signed [31:0] operation_194_3460;
wire [7:0] operation_194_3461;
reg signed [31:0] operation_194_3462;
wire [7:0] operation_194_3463;
reg signed [31:0] operation_194_3464;
wire [7:0] operation_194_3465;
reg signed [31:0] operation_194_3466;
wire [7:0] operation_194_3467;
reg signed [31:0] operation_194_3468;
wire [7:0] operation_194_3469;
reg signed [31:0] operation_194_3470;
wire [7:0] operation_194_3471;
reg signed [31:0] operation_194_3472;
wire [7:0] operation_194_3473;
reg signed [31:0] operation_194_3474;
wire [7:0] operation_194_3475;
reg signed [31:0] operation_194_3476;
wire signed [31:0] operation_194_3477;
wire signed [31:0] operation_194_3478;
wire signed [31:0] operation_194_3479;
wire signed [31:0] operation_194_3480;
wire signed [31:0] operation_194_3481;
wire signed [31:0] operation_194_3482;
wire signed [31:0] operation_194_3483;
wire signed [31:0] operation_194_3484;
wire signed [31:0] operation_194_3485;
wire signed [31:0] operation_194_3486;
wire signed [31:0] operation_194_3487;
wire signed [31:0] operation_194_3488;
wire signed [31:0] operation_194_3489;
wire signed [31:0] operation_194_3490;
wire signed [31:0] operation_194_3491;
wire signed [31:0] operation_194_3492;
wire signed [31:0] operation_194_3493;
wire signed [31:0] operation_194_3494;
wire [7:0] operation_194_3495;
reg signed [31:0] operation_194_3496;
wire [7:0] operation_194_3497;
reg signed [31:0] operation_194_3498;
wire [7:0] operation_194_3499;
reg signed [31:0] operation_194_3500;
wire [7:0] operation_194_3501;
reg signed [31:0] operation_194_3502;
wire [7:0] operation_194_3503;
reg signed [31:0] operation_194_3504;
wire [7:0] operation_194_3505;
reg signed [31:0] operation_194_3506;
wire [7:0] operation_194_3507;
reg signed [31:0] operation_194_3508;
wire [7:0] operation_194_3509;
reg signed [31:0] operation_194_3510;
wire [7:0] operation_194_3511;
reg signed [31:0] operation_194_3512;
wire [7:0] operation_194_3513;
reg signed [31:0] operation_194_3514;
wire signed [31:0] operation_194_3515;
wire signed [31:0] operation_194_3516;
wire signed [31:0] operation_194_3517;
wire signed [31:0] operation_194_3518;
wire signed [31:0] operation_194_3519;
wire signed [31:0] operation_194_3520;
wire signed [31:0] operation_194_3521;
wire signed [31:0] operation_194_3522;
wire signed [31:0] operation_194_3523;
wire signed [31:0] operation_194_3524;
wire [7:0] operation_194_3525;
reg signed [31:0] operation_194_3526;
wire [7:0] operation_194_3527;
reg signed [31:0] operation_194_3528;
wire [7:0] operation_194_3529;
reg signed [31:0] operation_194_3530;
wire [7:0] operation_194_3531;
reg signed [31:0] operation_194_3532;
wire [7:0] operation_194_3533;
reg signed [31:0] operation_194_3534;
wire [7:0] operation_194_3535;
reg signed [31:0] operation_194_3536;
wire [7:0] operation_194_3537;
reg signed [31:0] operation_194_3538;
wire [7:0] operation_194_3539;
reg signed [31:0] operation_194_3540;
wire [7:0] operation_194_3541;
reg signed [31:0] operation_194_3542;
wire [7:0] operation_194_3543;
reg signed [31:0] operation_194_3544;
wire signed [31:0] operation_194_3545;
wire signed [31:0] operation_194_3546;
wire signed [31:0] operation_194_3547;
wire signed [31:0] operation_194_3548;
wire signed [31:0] operation_194_3549;
wire signed [31:0] operation_194_3550;
wire signed [31:0] operation_194_3551;
wire signed [31:0] operation_194_3552;
wire signed [31:0] operation_194_3553;
wire signed [31:0] operation_194_3554;
wire [7:0] operation_194_3555;
reg signed [31:0] operation_194_3556;
wire [7:0] operation_194_3557;
reg signed [31:0] operation_194_3558;
wire [7:0] operation_194_3559;
reg signed [31:0] operation_194_3560;
wire [7:0] operation_194_3561;
reg signed [31:0] operation_194_3562;
wire [7:0] operation_194_3563;
reg signed [31:0] operation_194_3564;
wire [7:0] operation_194_3565;
reg signed [31:0] operation_194_3566;
wire [7:0] operation_194_3567;
reg signed [31:0] operation_194_3568;
wire [7:0] operation_194_3569;
reg signed [31:0] operation_194_3570;
wire [7:0] operation_194_3571;
reg signed [31:0] operation_194_3572;
wire [7:0] operation_194_3573;
reg signed [31:0] operation_194_3574;
wire signed [31:0] operation_194_3575;
wire signed [31:0] operation_194_3576;
wire signed [31:0] operation_194_3577;
wire signed [31:0] operation_194_3578;
wire signed [31:0] operation_194_3579;
wire signed [31:0] operation_194_3580;
wire signed [31:0] operation_194_3581;
wire signed [31:0] operation_194_3582;
wire signed [31:0] operation_194_3583;
wire signed [31:0] operation_194_3584;
wire [7:0] operation_194_3585;
reg signed [31:0] operation_194_3586;
reg signed [31:0] operation_194_3587;
wire [7:0] operation_194_3588;
reg signed [31:0] operation_194_3589;
reg signed [31:0] operation_194_3590;
wire [7:0] operation_194_3591;
reg signed [31:0] operation_194_3592;
reg signed [31:0] operation_194_3593;
wire [7:0] operation_194_3594;
reg signed [31:0] operation_194_3595;
reg signed [31:0] operation_194_3596;
wire [7:0] operation_194_3597;
reg signed [31:0] operation_194_3598;
reg signed [31:0] operation_194_3599;
wire [7:0] operation_194_3600;
reg signed [31:0] operation_194_3601;
reg signed [31:0] operation_194_3602;
wire [7:0] operation_194_3603;
reg signed [31:0] operation_194_3604;
reg signed [31:0] operation_194_3605;
wire [7:0] operation_194_3606;
reg signed [31:0] operation_194_3607;
reg signed [31:0] operation_194_3608;
wire [7:0] operation_194_3609;
reg signed [31:0] operation_194_3610;
wire [7:0] operation_194_3611;
reg signed [31:0] operation_194_3612;
wire signed [31:0] operation_194_3613;
wire signed [31:0] operation_194_3614;
reg signed [31:0] operation_194_3615;
reg signed [31:0] operation_194_3616;
reg signed [31:0] operation_194_3617;
wire signed [31:0] operation_194_3618;
reg signed [31:0] operation_194_3619;
reg signed [31:0] operation_194_3620;
reg signed [31:0] operation_194_3621;
wire signed [31:0] operation_194_3622;
reg signed [31:0] operation_194_3623;
reg signed [31:0] operation_194_3624;
reg signed [31:0] operation_194_3625;
wire signed [31:0] operation_194_3626;
reg signed [31:0] operation_194_3627;
reg signed [31:0] operation_194_3628;
reg signed [31:0] operation_194_3629;
wire signed [31:0] operation_194_3630;
reg signed [31:0] operation_194_3631;
reg signed [31:0] operation_194_3632;
reg signed [31:0] operation_194_3633;
wire signed [31:0] operation_194_3634;
reg signed [31:0] operation_194_3635;
reg signed [31:0] operation_194_3636;
reg signed [31:0] operation_194_3637;
wire signed [31:0] operation_194_3638;
reg signed [31:0] operation_194_3639;
reg signed [31:0] operation_194_3640;
reg signed [31:0] operation_194_3641;
wire signed [31:0] operation_194_3642;
reg signed [31:0] operation_194_3643;
reg signed [31:0] operation_194_3644;
reg signed [31:0] operation_194_3645;
wire signed [31:0] operation_194_3646;
wire [7:0] operation_194_3647;
reg signed [31:0] operation_194_3648;
reg signed [31:0] operation_194_3649;
wire [7:0] operation_194_3650;
reg signed [31:0] operation_194_3651;
reg signed [31:0] operation_194_3652;
wire [7:0] operation_194_3653;
reg signed [31:0] operation_194_3654;
reg signed [31:0] operation_194_3655;
wire [7:0] operation_194_3656;
reg signed [31:0] operation_194_3657;
reg signed [31:0] operation_194_3658;
wire [7:0] operation_194_3659;
reg signed [31:0] operation_194_3660;
reg signed [31:0] operation_194_3661;
wire [7:0] operation_194_3662;
reg signed [31:0] operation_194_3663;
reg signed [31:0] operation_194_3664;
wire [7:0] operation_194_3665;
reg signed [31:0] operation_194_3666;
reg signed [31:0] operation_194_3667;
wire [7:0] operation_194_3668;
reg signed [31:0] operation_194_3669;
reg signed [31:0] operation_194_3670;
wire [7:0] operation_194_3671;
reg signed [31:0] operation_194_3672;
wire [7:0] operation_194_3673;
reg signed [31:0] operation_194_3674;
wire signed [31:0] operation_194_3675;
wire signed [31:0] operation_194_3676;
wire signed [31:0] operation_194_3677;
wire signed [31:0] operation_194_3678;
reg signed [31:0] operation_194_3679;
reg signed [31:0] operation_194_3680;
reg signed [31:0] operation_194_3681;
wire signed [31:0] operation_194_3682;
reg signed [31:0] operation_194_3683;
reg signed [31:0] operation_194_3684;
reg signed [31:0] operation_194_3685;
wire signed [31:0] operation_194_3686;
reg signed [31:0] operation_194_3687;
reg signed [31:0] operation_194_3688;
reg signed [31:0] operation_194_3689;
wire signed [31:0] operation_194_3690;
reg signed [31:0] operation_194_3691;
reg signed [31:0] operation_194_3692;
reg signed [31:0] operation_194_3693;
wire signed [31:0] operation_194_3694;
reg signed [31:0] operation_194_3695;
reg signed [31:0] operation_194_3696;
reg signed [31:0] operation_194_3697;
wire signed [31:0] operation_194_3698;
reg signed [31:0] operation_194_3699;
reg signed [31:0] operation_194_3700;
reg signed [31:0] operation_194_3701;
wire signed [31:0] operation_194_3702;
reg signed [31:0] operation_194_3703;
reg signed [31:0] operation_194_3704;
reg signed [31:0] operation_194_3705;
wire signed [31:0] operation_194_3706;
reg signed [31:0] operation_194_3707;
reg signed [31:0] operation_194_3708;
reg signed [31:0] operation_194_3709;
wire signed [31:0] operation_194_3710;
wire [7:0] operation_194_3711;
wire [7:0] operation_194_3712;
reg signed [31:0] operation_194_3713;
wire [7:0] operation_194_3714;
wire [7:0] operation_194_3715;
reg signed [31:0] operation_194_3716;
wire [7:0] operation_194_3717;
wire [7:0] operation_194_3718;
reg signed [31:0] operation_194_3719;
wire [7:0] operation_194_3720;
wire [7:0] operation_194_3721;
reg signed [31:0] operation_194_3722;
wire [7:0] operation_194_3723;
reg signed [31:0] operation_194_3724;
wire [7:0] operation_194_3725;
reg signed [31:0] operation_194_3726;
wire [7:0] operation_194_3727;
reg signed [31:0] operation_194_3728;
wire [7:0] operation_194_3729;
reg signed [31:0] operation_194_3730;
wire [7:0] operation_194_3731;
reg signed [31:0] operation_194_3732;
wire signed [31:0] operation_194_3733;
wire signed [31:0] operation_194_3734;
wire signed [31:0] operation_194_3735;
wire signed [31:0] operation_194_3736;
wire signed [31:0] operation_194_3737;
reg signed [31:0] operation_194_3738;
reg signed [31:0] operation_194_3739;
reg signed [31:0] operation_194_3740;
reg signed [31:0] operation_194_3741;
wire [7:0] operation_194_3742;
reg signed [31:0] operation_194_3743;
wire [7:0] operation_194_3744;
reg signed [31:0] operation_194_3745;
wire [7:0] operation_194_3746;
reg signed [31:0] operation_194_3747;
wire [7:0] operation_194_3748;
reg signed [31:0] operation_194_3749;
wire [7:0] operation_194_3750;
reg signed [31:0] operation_194_3751;
wire [7:0] operation_194_3752;
reg signed [31:0] operation_194_3753;
wire [7:0] operation_194_3754;
reg signed [31:0] operation_194_3755;
wire [7:0] operation_194_3756;
reg signed [31:0] operation_194_3757;
wire [7:0] operation_194_3758;
reg signed [31:0] operation_194_3759;
wire [7:0] operation_194_3760;
reg signed [31:0] operation_194_3761;
wire [7:0] operation_194_3762;
reg signed [31:0] operation_194_3763;
wire signed [31:0] operation_194_3770;
reg signed [31:0] operation_194_3773;
reg signed [31:0] operation_194_3774;
reg signed [31:0] operation_194_3775;
reg signed [31:0] operation_194_3776;
wire signed [31:0] operation_194_3777;
wire signed [31:0] operation_194_3778;
wire signed [31:0] operation_194_3779;
wire signed [31:0] operation_194_3780;
wire signed [31:0] operation_194_3781;
wire signed [31:0] operation_194_3782;
wire signed [31:0] operation_194_3783;
wire signed [31:0] operation_194_3784;
wire [7:0] operation_194_3787;
reg signed [31:0] operation_194_3788;
wire [7:0] operation_194_3789;
reg signed [31:0] operation_194_3790;
wire signed [31:0] operation_194_3801;
wire signed [31:0] operation_194_3803;
reg [7:0] operation_194_3805_latch;
wire [7:0] operation_194_3805;
reg [7:0] operation_194_3806_latch;
wire [7:0] operation_194_3806;
wire signed [31:0] operation_194_3807;
wire signed [31:0] operation_194_3808;
wire signed [31:0] operation_194_3809;
wire signed [31:0] operation_194_3810;
wire signed [31:0] operation_194_3811;
wire signed [31:0] operation_194_3812;
wire signed [31:0] operation_194_3813;
wire signed [31:0] operation_194_3814;
reg [7:0] operation_194_3815_latch;
wire [7:0] operation_194_3815;
reg [7:0] operation_194_3816_latch;
wire [7:0] operation_194_3816;
reg [7:0] operation_194_3817_latch;
wire [7:0] operation_194_3817;
reg [7:0] operation_194_3818_latch;
wire [7:0] operation_194_3818;
reg [7:0] operation_194_3819_latch;
wire [7:0] operation_194_3819;
reg [7:0] operation_194_3820_latch;
wire [7:0] operation_194_3820;
reg [7:0] operation_194_3821_latch;
wire [7:0] operation_194_3821;
reg [7:0] operation_194_3822_latch;
wire [7:0] operation_194_3822;
reg [7:0] operation_194_3823_latch;
wire [7:0] operation_194_3823;
reg [7:0] operation_194_3824_latch;
wire [7:0] operation_194_3824;
reg [7:0] operation_194_3825_latch;
wire [7:0] operation_194_3825;
reg [7:0] operation_194_3826_latch;
wire [7:0] operation_194_3826;
reg [7:0] operation_194_3827_latch;
wire [7:0] operation_194_3827;
reg [7:0] operation_194_3828_latch;
wire [7:0] operation_194_3828;
reg [7:0] operation_194_3829_latch;
wire [7:0] operation_194_3829;
reg [7:0] operation_194_3830_latch;
wire [7:0] operation_194_3830;
reg [7:0] operation_194_3831_latch;
wire [7:0] operation_194_3831;
reg [7:0] operation_194_3832_latch;
wire [7:0] operation_194_3832;
wire [7:0] operation_194_2986;
reg signed [31:0] operation_194_2987;
wire signed [31:0] operation_194_2988;
wire [7:0] operation_194_2990;
reg signed [31:0] operation_194_2991;
wire [7:0] operation_194_2992;
reg signed [31:0] operation_194_2993;
wire [7:0] operation_194_2994;
reg signed [31:0] operation_194_2995;
wire [7:0] operation_194_2996;
reg signed [31:0] operation_194_2997;
wire [7:0] operation_194_2998;
reg signed [31:0] operation_194_2999;
wire [7:0] operation_194_3000;
reg signed [31:0] operation_194_3001;
wire [7:0] operation_194_3002;
reg signed [31:0] operation_194_3003;
wire [7:0] operation_194_3004;
reg signed [31:0] operation_194_3005;
wire signed [31:0] operation_194_3006;
wire signed [31:0] operation_194_3007;
wire signed [31:0] operation_194_3008;
wire signed [31:0] operation_194_3009;
wire signed [31:0] operation_194_3010;
wire signed [31:0] operation_194_3011;
wire signed [31:0] operation_194_3012;
wire signed [31:0] operation_194_3013;
wire signed [31:0] operation_194_3014;
wire signed [31:0] operation_194_3015;
wire [7:0] operation_194_3016;
reg signed [31:0] operation_194_3017;
wire [7:0] operation_194_3018;
reg signed [31:0] operation_194_3019;
wire [7:0] operation_194_3020;
reg signed [31:0] operation_194_3021;
wire [7:0] operation_194_3022;
reg signed [31:0] operation_194_3023;
wire [7:0] operation_194_3024;
reg signed [31:0] operation_194_3025;
wire [7:0] operation_194_3026;
reg signed [31:0] operation_194_3027;
wire [7:0] operation_194_3028;
reg signed [31:0] operation_194_3029;
wire [7:0] operation_194_3030;
reg signed [31:0] operation_194_3031;
wire [7:0] operation_194_3032;
reg signed [31:0] operation_194_3033;
wire [7:0] operation_194_3034;
reg signed [31:0] operation_194_3035;
wire [7:0] operation_194_3036;
reg signed [31:0] operation_194_3037;
wire [7:0] operation_194_3038;
reg signed [31:0] operation_194_3039;
wire [7:0] operation_194_3040;
reg signed [31:0] operation_194_3041;
wire [7:0] operation_194_3042;
reg signed [31:0] operation_194_3043;
wire [7:0] operation_194_3044;
reg signed [31:0] operation_194_3045;
wire [7:0] operation_194_3046;
reg signed [31:0] operation_194_3047;
wire signed [31:0] operation_194_3048;
wire signed [31:0] operation_194_3049;
wire signed [31:0] operation_194_3050;
wire signed [31:0] operation_194_3051;
wire signed [31:0] operation_194_3052;
wire signed [31:0] operation_194_3053;
wire signed [31:0] operation_194_3054;
wire signed [31:0] operation_194_3055;
wire signed [31:0] operation_194_3056;
wire signed [31:0] operation_194_3057;
wire signed [31:0] operation_194_3058;
wire signed [31:0] operation_194_3059;
wire signed [31:0] operation_194_3060;
wire signed [31:0] operation_194_3061;
wire signed [31:0] operation_194_3062;
wire signed [31:0] operation_194_3063;
wire signed [31:0] operation_194_3064;
wire signed [31:0] operation_194_3065;
wire [7:0] operation_194_3066;
reg signed [31:0] operation_194_3067;
wire [7:0] operation_194_3068;
reg signed [31:0] operation_194_3069;
wire [7:0] operation_194_3070;
reg signed [31:0] operation_194_3071;
wire [7:0] operation_194_3072;
reg signed [31:0] operation_194_3073;
wire [7:0] operation_194_3074;
reg signed [31:0] operation_194_3075;
wire [7:0] operation_194_3076;
reg signed [31:0] operation_194_3077;
wire [7:0] operation_194_3078;
reg signed [31:0] operation_194_3079;
wire [7:0] operation_194_3080;
reg signed [31:0] operation_194_3081;
wire [7:0] operation_194_3082;
reg signed [31:0] operation_194_3083;
wire [7:0] operation_194_3084;
reg signed [31:0] operation_194_3085;
wire signed [31:0] operation_194_3086;
wire signed [31:0] operation_194_3087;
wire signed [31:0] operation_194_3088;
wire signed [31:0] operation_194_3089;
wire signed [31:0] operation_194_3090;
wire signed [31:0] operation_194_3091;
wire signed [31:0] operation_194_3092;
wire signed [31:0] operation_194_3093;
wire signed [31:0] operation_194_3094;
wire signed [31:0] operation_194_3095;
wire [7:0] operation_194_3096;
reg signed [31:0] operation_194_3097;
wire [7:0] operation_194_3098;
reg signed [31:0] operation_194_3099;
wire [7:0] operation_194_3100;
reg signed [31:0] operation_194_3101;
wire [7:0] operation_194_3102;
reg signed [31:0] operation_194_3103;
wire [7:0] operation_194_3104;
reg signed [31:0] operation_194_3105;
wire [7:0] operation_194_3106;
reg signed [31:0] operation_194_3107;
wire [7:0] operation_194_3108;
reg signed [31:0] operation_194_3109;
wire [7:0] operation_194_3110;
reg signed [31:0] operation_194_3111;
wire [7:0] operation_194_3112;
reg signed [31:0] operation_194_3113;
wire [7:0] operation_194_3114;
reg signed [31:0] operation_194_3115;
wire signed [31:0] operation_194_3116;
wire signed [31:0] operation_194_3117;
wire signed [31:0] operation_194_3118;
wire signed [31:0] operation_194_3119;
wire signed [31:0] operation_194_3120;
wire signed [31:0] operation_194_3121;
wire signed [31:0] operation_194_3122;
wire signed [31:0] operation_194_3123;
wire signed [31:0] operation_194_3124;
wire signed [31:0] operation_194_3125;
wire [7:0] operation_194_3126;
reg signed [31:0] operation_194_3127;
wire [7:0] operation_194_3128;
reg signed [31:0] operation_194_3129;
wire [7:0] operation_194_3130;
reg signed [31:0] operation_194_3131;
wire [7:0] operation_194_3132;
reg signed [31:0] operation_194_3133;
wire [7:0] operation_194_3134;
reg signed [31:0] operation_194_3135;
wire [7:0] operation_194_3136;
reg signed [31:0] operation_194_3137;
wire [7:0] operation_194_3138;
reg signed [31:0] operation_194_3139;
wire [7:0] operation_194_3140;
reg signed [31:0] operation_194_3141;
wire [7:0] operation_194_3142;
reg signed [31:0] operation_194_3143;
wire [7:0] operation_194_3144;
reg signed [31:0] operation_194_3145;
wire signed [31:0] operation_194_3146;
wire signed [31:0] operation_194_3147;
wire signed [31:0] operation_194_3148;
wire signed [31:0] operation_194_3149;
wire signed [31:0] operation_194_3150;
wire signed [31:0] operation_194_3151;
wire signed [31:0] operation_194_3152;
wire signed [31:0] operation_194_3153;
wire signed [31:0] operation_194_3154;
wire signed [31:0] operation_194_3155;
wire [7:0] operation_194_3156;
reg signed [31:0] operation_194_3157;
reg signed [31:0] operation_194_3158;
wire [7:0] operation_194_3159;
reg signed [31:0] operation_194_3160;
reg signed [31:0] operation_194_3161;
wire [7:0] operation_194_3162;
reg signed [31:0] operation_194_3163;
reg signed [31:0] operation_194_3164;
wire [7:0] operation_194_3165;
reg signed [31:0] operation_194_3166;
reg signed [31:0] operation_194_3167;
wire [7:0] operation_194_3168;
reg signed [31:0] operation_194_3169;
reg signed [31:0] operation_194_3170;
wire [7:0] operation_194_3171;
reg signed [31:0] operation_194_3172;
reg signed [31:0] operation_194_3173;
wire [7:0] operation_194_3174;
reg signed [31:0] operation_194_3175;
reg signed [31:0] operation_194_3176;
wire [7:0] operation_194_3177;
reg signed [31:0] operation_194_3178;
reg signed [31:0] operation_194_3179;
wire [7:0] operation_194_3180;
reg signed [31:0] operation_194_3181;
wire [7:0] operation_194_3182;
reg signed [31:0] operation_194_3183;
wire signed [31:0] operation_194_3184;
wire signed [31:0] operation_194_3185;
reg signed [31:0] operation_194_3186;
reg signed [31:0] operation_194_3187;
reg signed [31:0] operation_194_3188;
wire signed [31:0] operation_194_3189;
reg signed [31:0] operation_194_3190;
reg signed [31:0] operation_194_3191;
reg signed [31:0] operation_194_3192;
wire signed [31:0] operation_194_3193;
reg signed [31:0] operation_194_3194;
reg signed [31:0] operation_194_3195;
reg signed [31:0] operation_194_3196;
wire signed [31:0] operation_194_3197;
reg signed [31:0] operation_194_3198;
reg signed [31:0] operation_194_3199;
reg signed [31:0] operation_194_3200;
wire signed [31:0] operation_194_3201;
reg signed [31:0] operation_194_3202;
reg signed [31:0] operation_194_3203;
reg signed [31:0] operation_194_3204;
wire signed [31:0] operation_194_3205;
reg signed [31:0] operation_194_3206;
reg signed [31:0] operation_194_3207;
reg signed [31:0] operation_194_3208;
wire signed [31:0] operation_194_3209;
reg signed [31:0] operation_194_3210;
reg signed [31:0] operation_194_3211;
reg signed [31:0] operation_194_3212;
wire signed [31:0] operation_194_3213;
reg signed [31:0] operation_194_3214;
reg signed [31:0] operation_194_3215;
reg signed [31:0] operation_194_3216;
wire signed [31:0] operation_194_3217;
wire [7:0] operation_194_3218;
reg signed [31:0] operation_194_3219;
reg signed [31:0] operation_194_3220;
wire [7:0] operation_194_3221;
reg signed [31:0] operation_194_3222;
reg signed [31:0] operation_194_3223;
wire [7:0] operation_194_3224;
reg signed [31:0] operation_194_3225;
reg signed [31:0] operation_194_3226;
wire [7:0] operation_194_3227;
reg signed [31:0] operation_194_3228;
reg signed [31:0] operation_194_3229;
wire [7:0] operation_194_3230;
reg signed [31:0] operation_194_3231;
reg signed [31:0] operation_194_3232;
wire [7:0] operation_194_3233;
reg signed [31:0] operation_194_3234;
reg signed [31:0] operation_194_3235;
wire [7:0] operation_194_3236;
reg signed [31:0] operation_194_3237;
reg signed [31:0] operation_194_3238;
wire [7:0] operation_194_3239;
reg signed [31:0] operation_194_3240;
reg signed [31:0] operation_194_3241;
wire [7:0] operation_194_3242;
reg signed [31:0] operation_194_3243;
wire [7:0] operation_194_3244;
reg signed [31:0] operation_194_3245;
wire signed [31:0] operation_194_3246;
wire signed [31:0] operation_194_3247;
wire signed [31:0] operation_194_3248;
wire signed [31:0] operation_194_3249;
reg signed [31:0] operation_194_3250;
reg signed [31:0] operation_194_3251;
reg signed [31:0] operation_194_3252;
wire signed [31:0] operation_194_3253;
reg signed [31:0] operation_194_3254;
reg signed [31:0] operation_194_3255;
reg signed [31:0] operation_194_3256;
wire signed [31:0] operation_194_3257;
reg signed [31:0] operation_194_3258;
reg signed [31:0] operation_194_3259;
reg signed [31:0] operation_194_3260;
wire signed [31:0] operation_194_3261;
reg signed [31:0] operation_194_3262;
reg signed [31:0] operation_194_3263;
reg signed [31:0] operation_194_3264;
wire signed [31:0] operation_194_3265;
reg signed [31:0] operation_194_3266;
reg signed [31:0] operation_194_3267;
reg signed [31:0] operation_194_3268;
wire signed [31:0] operation_194_3269;
reg signed [31:0] operation_194_3270;
reg signed [31:0] operation_194_3271;
reg signed [31:0] operation_194_3272;
wire signed [31:0] operation_194_3273;
reg signed [31:0] operation_194_3274;
reg signed [31:0] operation_194_3275;
reg signed [31:0] operation_194_3276;
wire signed [31:0] operation_194_3277;
reg signed [31:0] operation_194_3278;
reg signed [31:0] operation_194_3279;
reg signed [31:0] operation_194_3280;
wire signed [31:0] operation_194_3281;
wire [7:0] operation_194_3282;
wire [7:0] operation_194_3283;
reg signed [31:0] operation_194_3284;
wire [7:0] operation_194_3285;
wire [7:0] operation_194_3286;
reg signed [31:0] operation_194_3287;
wire [7:0] operation_194_3288;
wire [7:0] operation_194_3289;
reg signed [31:0] operation_194_3290;
wire [7:0] operation_194_3291;
wire [7:0] operation_194_3292;
reg signed [31:0] operation_194_3293;
wire [7:0] operation_194_3294;
reg signed [31:0] operation_194_3295;
wire [7:0] operation_194_3296;
reg signed [31:0] operation_194_3297;
wire [7:0] operation_194_3298;
reg signed [31:0] operation_194_3299;
wire [7:0] operation_194_3300;
reg signed [31:0] operation_194_3301;
wire [7:0] operation_194_3302;
reg signed [31:0] operation_194_3303;
wire signed [31:0] operation_194_3304;
wire signed [31:0] operation_194_3305;
wire signed [31:0] operation_194_3306;
wire signed [31:0] operation_194_3307;
wire signed [31:0] operation_194_3308;
reg signed [31:0] operation_194_3309;
reg signed [31:0] operation_194_3310;
reg signed [31:0] operation_194_3311;
reg signed [31:0] operation_194_3312;
wire [7:0] operation_194_3313;
reg signed [31:0] operation_194_3314;
wire [7:0] operation_194_3315;
reg signed [31:0] operation_194_3316;
wire [7:0] operation_194_3317;
reg signed [31:0] operation_194_3318;
wire [7:0] operation_194_3319;
reg signed [31:0] operation_194_3320;
wire [7:0] operation_194_3321;
reg signed [31:0] operation_194_3322;
wire [7:0] operation_194_3323;
reg signed [31:0] operation_194_3324;
wire [7:0] operation_194_3325;
reg signed [31:0] operation_194_3326;
wire [7:0] operation_194_3327;
reg signed [31:0] operation_194_3328;
wire [7:0] operation_194_3329;
reg signed [31:0] operation_194_3330;
wire [7:0] operation_194_3331;
reg signed [31:0] operation_194_3332;
wire [7:0] operation_194_3333;
reg signed [31:0] operation_194_3334;
wire signed [31:0] operation_194_3341;
reg signed [31:0] operation_194_3344;
reg signed [31:0] operation_194_3345;
reg signed [31:0] operation_194_3346;
reg signed [31:0] operation_194_3347;
wire signed [31:0] operation_194_3348;
wire signed [31:0] operation_194_3349;
wire signed [31:0] operation_194_3350;
wire signed [31:0] operation_194_3351;
wire signed [31:0] operation_194_3352;
wire signed [31:0] operation_194_3353;
wire signed [31:0] operation_194_3354;
wire signed [31:0] operation_194_3355;
wire [7:0] operation_194_3358;
reg signed [31:0] operation_194_3359;
wire [7:0] operation_194_3360;
reg signed [31:0] operation_194_3361;
wire signed [31:0] operation_194_3372;
wire signed [31:0] operation_194_3374;
reg [7:0] operation_194_3376_latch;
wire [7:0] operation_194_3376;
reg [7:0] operation_194_3377_latch;
wire [7:0] operation_194_3377;
wire signed [31:0] operation_194_3378;
wire signed [31:0] operation_194_3379;
wire signed [31:0] operation_194_3380;
wire signed [31:0] operation_194_3381;
wire signed [31:0] operation_194_3382;
wire signed [31:0] operation_194_3383;
wire signed [31:0] operation_194_3384;
wire signed [31:0] operation_194_3385;
reg [7:0] operation_194_3386_latch;
wire [7:0] operation_194_3386;
reg [7:0] operation_194_3387_latch;
wire [7:0] operation_194_3387;
reg [7:0] operation_194_3388_latch;
wire [7:0] operation_194_3388;
reg [7:0] operation_194_3389_latch;
wire [7:0] operation_194_3389;
reg [7:0] operation_194_3390_latch;
wire [7:0] operation_194_3390;
reg [7:0] operation_194_3391_latch;
wire [7:0] operation_194_3391;
reg [7:0] operation_194_3392_latch;
wire [7:0] operation_194_3392;
reg [7:0] operation_194_3393_latch;
wire [7:0] operation_194_3393;
reg [7:0] operation_194_3394_latch;
wire [7:0] operation_194_3394;
reg [7:0] operation_194_3395_latch;
wire [7:0] operation_194_3395;
reg [7:0] operation_194_3396_latch;
wire [7:0] operation_194_3396;
reg [7:0] operation_194_3397_latch;
wire [7:0] operation_194_3397;
reg [7:0] operation_194_3398_latch;
wire [7:0] operation_194_3398;
reg [7:0] operation_194_3399_latch;
wire [7:0] operation_194_3399;
reg [7:0] operation_194_3400_latch;
wire [7:0] operation_194_3400;
reg [7:0] operation_194_3401_latch;
wire [7:0] operation_194_3401;
reg [7:0] operation_194_3402_latch;
wire [7:0] operation_194_3402;
reg [7:0] operation_194_3403_latch;
wire [7:0] operation_194_3403;
wire [7:0] operation_194_2557;
reg signed [31:0] operation_194_2558;
wire signed [31:0] operation_194_2559;
wire [7:0] operation_194_2561;
reg signed [31:0] operation_194_2562;
wire [7:0] operation_194_2563;
reg signed [31:0] operation_194_2564;
wire [7:0] operation_194_2565;
reg signed [31:0] operation_194_2566;
wire [7:0] operation_194_2567;
reg signed [31:0] operation_194_2568;
wire [7:0] operation_194_2569;
reg signed [31:0] operation_194_2570;
wire [7:0] operation_194_2571;
reg signed [31:0] operation_194_2572;
wire [7:0] operation_194_2573;
reg signed [31:0] operation_194_2574;
wire [7:0] operation_194_2575;
reg signed [31:0] operation_194_2576;
wire signed [31:0] operation_194_2577;
wire signed [31:0] operation_194_2578;
wire signed [31:0] operation_194_2579;
wire signed [31:0] operation_194_2580;
wire signed [31:0] operation_194_2581;
wire signed [31:0] operation_194_2582;
wire signed [31:0] operation_194_2583;
wire signed [31:0] operation_194_2584;
wire signed [31:0] operation_194_2585;
wire signed [31:0] operation_194_2586;
wire [7:0] operation_194_2587;
reg signed [31:0] operation_194_2588;
wire [7:0] operation_194_2589;
reg signed [31:0] operation_194_2590;
wire [7:0] operation_194_2591;
reg signed [31:0] operation_194_2592;
wire [7:0] operation_194_2593;
reg signed [31:0] operation_194_2594;
wire [7:0] operation_194_2595;
reg signed [31:0] operation_194_2596;
wire [7:0] operation_194_2597;
reg signed [31:0] operation_194_2598;
wire [7:0] operation_194_2599;
reg signed [31:0] operation_194_2600;
wire [7:0] operation_194_2601;
reg signed [31:0] operation_194_2602;
wire [7:0] operation_194_2603;
reg signed [31:0] operation_194_2604;
wire [7:0] operation_194_2605;
reg signed [31:0] operation_194_2606;
wire [7:0] operation_194_2607;
reg signed [31:0] operation_194_2608;
wire [7:0] operation_194_2609;
reg signed [31:0] operation_194_2610;
wire [7:0] operation_194_2611;
reg signed [31:0] operation_194_2612;
wire [7:0] operation_194_2613;
reg signed [31:0] operation_194_2614;
wire [7:0] operation_194_2615;
reg signed [31:0] operation_194_2616;
wire [7:0] operation_194_2617;
reg signed [31:0] operation_194_2618;
wire signed [31:0] operation_194_2619;
wire signed [31:0] operation_194_2620;
wire signed [31:0] operation_194_2621;
wire signed [31:0] operation_194_2622;
wire signed [31:0] operation_194_2623;
wire signed [31:0] operation_194_2624;
wire signed [31:0] operation_194_2625;
wire signed [31:0] operation_194_2626;
wire signed [31:0] operation_194_2627;
wire signed [31:0] operation_194_2628;
wire signed [31:0] operation_194_2629;
wire signed [31:0] operation_194_2630;
wire signed [31:0] operation_194_2631;
wire signed [31:0] operation_194_2632;
wire signed [31:0] operation_194_2633;
wire signed [31:0] operation_194_2634;
wire signed [31:0] operation_194_2635;
wire signed [31:0] operation_194_2636;
wire [7:0] operation_194_2637;
reg signed [31:0] operation_194_2638;
wire [7:0] operation_194_2639;
reg signed [31:0] operation_194_2640;
wire [7:0] operation_194_2641;
reg signed [31:0] operation_194_2642;
wire [7:0] operation_194_2643;
reg signed [31:0] operation_194_2644;
wire [7:0] operation_194_2645;
reg signed [31:0] operation_194_2646;
wire [7:0] operation_194_2647;
reg signed [31:0] operation_194_2648;
wire [7:0] operation_194_2649;
reg signed [31:0] operation_194_2650;
wire [7:0] operation_194_2651;
reg signed [31:0] operation_194_2652;
wire [7:0] operation_194_2653;
reg signed [31:0] operation_194_2654;
wire [7:0] operation_194_2655;
reg signed [31:0] operation_194_2656;
wire signed [31:0] operation_194_2657;
wire signed [31:0] operation_194_2658;
wire signed [31:0] operation_194_2659;
wire signed [31:0] operation_194_2660;
wire signed [31:0] operation_194_2661;
wire signed [31:0] operation_194_2662;
wire signed [31:0] operation_194_2663;
wire signed [31:0] operation_194_2664;
wire signed [31:0] operation_194_2665;
wire signed [31:0] operation_194_2666;
wire [7:0] operation_194_2667;
reg signed [31:0] operation_194_2668;
wire [7:0] operation_194_2669;
reg signed [31:0] operation_194_2670;
wire [7:0] operation_194_2671;
reg signed [31:0] operation_194_2672;
wire [7:0] operation_194_2673;
reg signed [31:0] operation_194_2674;
wire [7:0] operation_194_2675;
reg signed [31:0] operation_194_2676;
wire [7:0] operation_194_2677;
reg signed [31:0] operation_194_2678;
wire [7:0] operation_194_2679;
reg signed [31:0] operation_194_2680;
wire [7:0] operation_194_2681;
reg signed [31:0] operation_194_2682;
wire [7:0] operation_194_2683;
reg signed [31:0] operation_194_2684;
wire [7:0] operation_194_2685;
reg signed [31:0] operation_194_2686;
wire signed [31:0] operation_194_2687;
wire signed [31:0] operation_194_2688;
wire signed [31:0] operation_194_2689;
wire signed [31:0] operation_194_2690;
wire signed [31:0] operation_194_2691;
wire signed [31:0] operation_194_2692;
wire signed [31:0] operation_194_2693;
wire signed [31:0] operation_194_2694;
wire signed [31:0] operation_194_2695;
wire signed [31:0] operation_194_2696;
wire [7:0] operation_194_2697;
reg signed [31:0] operation_194_2698;
wire [7:0] operation_194_2699;
reg signed [31:0] operation_194_2700;
wire [7:0] operation_194_2701;
reg signed [31:0] operation_194_2702;
wire [7:0] operation_194_2703;
reg signed [31:0] operation_194_2704;
wire [7:0] operation_194_2705;
reg signed [31:0] operation_194_2706;
wire [7:0] operation_194_2707;
reg signed [31:0] operation_194_2708;
wire [7:0] operation_194_2709;
reg signed [31:0] operation_194_2710;
wire [7:0] operation_194_2711;
reg signed [31:0] operation_194_2712;
wire [7:0] operation_194_2713;
reg signed [31:0] operation_194_2714;
wire [7:0] operation_194_2715;
reg signed [31:0] operation_194_2716;
wire signed [31:0] operation_194_2717;
wire signed [31:0] operation_194_2718;
wire signed [31:0] operation_194_2719;
wire signed [31:0] operation_194_2720;
wire signed [31:0] operation_194_2721;
wire signed [31:0] operation_194_2722;
wire signed [31:0] operation_194_2723;
wire signed [31:0] operation_194_2724;
wire signed [31:0] operation_194_2725;
wire signed [31:0] operation_194_2726;
wire [7:0] operation_194_2727;
reg signed [31:0] operation_194_2728;
reg signed [31:0] operation_194_2729;
wire [7:0] operation_194_2730;
reg signed [31:0] operation_194_2731;
reg signed [31:0] operation_194_2732;
wire [7:0] operation_194_2733;
reg signed [31:0] operation_194_2734;
reg signed [31:0] operation_194_2735;
wire [7:0] operation_194_2736;
reg signed [31:0] operation_194_2737;
reg signed [31:0] operation_194_2738;
wire [7:0] operation_194_2739;
reg signed [31:0] operation_194_2740;
reg signed [31:0] operation_194_2741;
wire [7:0] operation_194_2742;
reg signed [31:0] operation_194_2743;
reg signed [31:0] operation_194_2744;
wire [7:0] operation_194_2745;
reg signed [31:0] operation_194_2746;
reg signed [31:0] operation_194_2747;
wire [7:0] operation_194_2748;
reg signed [31:0] operation_194_2749;
reg signed [31:0] operation_194_2750;
wire [7:0] operation_194_2751;
reg signed [31:0] operation_194_2752;
wire [7:0] operation_194_2753;
reg signed [31:0] operation_194_2754;
wire signed [31:0] operation_194_2755;
wire signed [31:0] operation_194_2756;
reg signed [31:0] operation_194_2757;
reg signed [31:0] operation_194_2758;
reg signed [31:0] operation_194_2759;
wire signed [31:0] operation_194_2760;
reg signed [31:0] operation_194_2761;
reg signed [31:0] operation_194_2762;
reg signed [31:0] operation_194_2763;
wire signed [31:0] operation_194_2764;
reg signed [31:0] operation_194_2765;
reg signed [31:0] operation_194_2766;
reg signed [31:0] operation_194_2767;
wire signed [31:0] operation_194_2768;
reg signed [31:0] operation_194_2769;
reg signed [31:0] operation_194_2770;
reg signed [31:0] operation_194_2771;
wire signed [31:0] operation_194_2772;
reg signed [31:0] operation_194_2773;
reg signed [31:0] operation_194_2774;
reg signed [31:0] operation_194_2775;
wire signed [31:0] operation_194_2776;
reg signed [31:0] operation_194_2777;
reg signed [31:0] operation_194_2778;
reg signed [31:0] operation_194_2779;
wire signed [31:0] operation_194_2780;
reg signed [31:0] operation_194_2781;
reg signed [31:0] operation_194_2782;
reg signed [31:0] operation_194_2783;
wire signed [31:0] operation_194_2784;
reg signed [31:0] operation_194_2785;
reg signed [31:0] operation_194_2786;
reg signed [31:0] operation_194_2787;
wire signed [31:0] operation_194_2788;
wire [7:0] operation_194_2789;
reg signed [31:0] operation_194_2790;
reg signed [31:0] operation_194_2791;
wire [7:0] operation_194_2792;
reg signed [31:0] operation_194_2793;
reg signed [31:0] operation_194_2794;
wire [7:0] operation_194_2795;
reg signed [31:0] operation_194_2796;
reg signed [31:0] operation_194_2797;
wire [7:0] operation_194_2798;
reg signed [31:0] operation_194_2799;
reg signed [31:0] operation_194_2800;
wire [7:0] operation_194_2801;
reg signed [31:0] operation_194_2802;
reg signed [31:0] operation_194_2803;
wire [7:0] operation_194_2804;
reg signed [31:0] operation_194_2805;
reg signed [31:0] operation_194_2806;
wire [7:0] operation_194_2807;
reg signed [31:0] operation_194_2808;
reg signed [31:0] operation_194_2809;
wire [7:0] operation_194_2810;
reg signed [31:0] operation_194_2811;
reg signed [31:0] operation_194_2812;
wire [7:0] operation_194_2813;
reg signed [31:0] operation_194_2814;
wire [7:0] operation_194_2815;
reg signed [31:0] operation_194_2816;
wire signed [31:0] operation_194_2817;
wire signed [31:0] operation_194_2818;
wire signed [31:0] operation_194_2819;
wire signed [31:0] operation_194_2820;
reg signed [31:0] operation_194_2821;
reg signed [31:0] operation_194_2822;
reg signed [31:0] operation_194_2823;
wire signed [31:0] operation_194_2824;
reg signed [31:0] operation_194_2825;
reg signed [31:0] operation_194_2826;
reg signed [31:0] operation_194_2827;
wire signed [31:0] operation_194_2828;
reg signed [31:0] operation_194_2829;
reg signed [31:0] operation_194_2830;
reg signed [31:0] operation_194_2831;
wire signed [31:0] operation_194_2832;
reg signed [31:0] operation_194_2833;
reg signed [31:0] operation_194_2834;
reg signed [31:0] operation_194_2835;
wire signed [31:0] operation_194_2836;
reg signed [31:0] operation_194_2837;
reg signed [31:0] operation_194_2838;
reg signed [31:0] operation_194_2839;
wire signed [31:0] operation_194_2840;
reg signed [31:0] operation_194_2841;
reg signed [31:0] operation_194_2842;
reg signed [31:0] operation_194_2843;
wire signed [31:0] operation_194_2844;
reg signed [31:0] operation_194_2845;
reg signed [31:0] operation_194_2846;
reg signed [31:0] operation_194_2847;
wire signed [31:0] operation_194_2848;
reg signed [31:0] operation_194_2849;
reg signed [31:0] operation_194_2850;
reg signed [31:0] operation_194_2851;
wire signed [31:0] operation_194_2852;
wire [7:0] operation_194_2853;
wire [7:0] operation_194_2854;
reg signed [31:0] operation_194_2855;
wire [7:0] operation_194_2856;
wire [7:0] operation_194_2857;
reg signed [31:0] operation_194_2858;
wire [7:0] operation_194_2859;
wire [7:0] operation_194_2860;
reg signed [31:0] operation_194_2861;
wire [7:0] operation_194_2862;
wire [7:0] operation_194_2863;
reg signed [31:0] operation_194_2864;
wire [7:0] operation_194_2865;
reg signed [31:0] operation_194_2866;
wire [7:0] operation_194_2867;
reg signed [31:0] operation_194_2868;
wire [7:0] operation_194_2869;
reg signed [31:0] operation_194_2870;
wire [7:0] operation_194_2871;
reg signed [31:0] operation_194_2872;
wire [7:0] operation_194_2873;
reg signed [31:0] operation_194_2874;
wire signed [31:0] operation_194_2875;
wire signed [31:0] operation_194_2876;
wire signed [31:0] operation_194_2877;
wire signed [31:0] operation_194_2878;
wire signed [31:0] operation_194_2879;
reg signed [31:0] operation_194_2880;
reg signed [31:0] operation_194_2881;
reg signed [31:0] operation_194_2882;
reg signed [31:0] operation_194_2883;
wire [7:0] operation_194_2884;
reg signed [31:0] operation_194_2885;
wire [7:0] operation_194_2886;
reg signed [31:0] operation_194_2887;
wire [7:0] operation_194_2888;
reg signed [31:0] operation_194_2889;
wire [7:0] operation_194_2890;
reg signed [31:0] operation_194_2891;
wire [7:0] operation_194_2892;
reg signed [31:0] operation_194_2893;
wire [7:0] operation_194_2894;
reg signed [31:0] operation_194_2895;
wire [7:0] operation_194_2896;
reg signed [31:0] operation_194_2897;
wire [7:0] operation_194_2898;
reg signed [31:0] operation_194_2899;
wire [7:0] operation_194_2900;
reg signed [31:0] operation_194_2901;
wire [7:0] operation_194_2902;
reg signed [31:0] operation_194_2903;
wire [7:0] operation_194_2904;
reg signed [31:0] operation_194_2905;
wire signed [31:0] operation_194_2912;
reg signed [31:0] operation_194_2915;
reg signed [31:0] operation_194_2916;
reg signed [31:0] operation_194_2917;
reg signed [31:0] operation_194_2918;
wire signed [31:0] operation_194_2919;
wire signed [31:0] operation_194_2920;
wire signed [31:0] operation_194_2921;
wire signed [31:0] operation_194_2922;
wire signed [31:0] operation_194_2923;
wire signed [31:0] operation_194_2924;
wire signed [31:0] operation_194_2925;
wire signed [31:0] operation_194_2926;
wire [7:0] operation_194_2929;
reg signed [31:0] operation_194_2930;
wire [7:0] operation_194_2931;
reg signed [31:0] operation_194_2932;
wire signed [31:0] operation_194_2943;
wire signed [31:0] operation_194_2945;
reg [7:0] operation_194_2947_latch;
wire [7:0] operation_194_2947;
reg [7:0] operation_194_2948_latch;
wire [7:0] operation_194_2948;
wire signed [31:0] operation_194_2949;
wire signed [31:0] operation_194_2950;
wire signed [31:0] operation_194_2951;
wire signed [31:0] operation_194_2952;
wire signed [31:0] operation_194_2953;
wire signed [31:0] operation_194_2954;
wire signed [31:0] operation_194_2955;
wire signed [31:0] operation_194_2956;
reg [7:0] operation_194_2957_latch;
wire [7:0] operation_194_2957;
reg [7:0] operation_194_2958_latch;
wire [7:0] operation_194_2958;
reg [7:0] operation_194_2959_latch;
wire [7:0] operation_194_2959;
reg [7:0] operation_194_2960_latch;
wire [7:0] operation_194_2960;
reg [7:0] operation_194_2961_latch;
wire [7:0] operation_194_2961;
reg [7:0] operation_194_2962_latch;
wire [7:0] operation_194_2962;
reg [7:0] operation_194_2963_latch;
wire [7:0] operation_194_2963;
reg [7:0] operation_194_2964_latch;
wire [7:0] operation_194_2964;
reg [7:0] operation_194_2965_latch;
wire [7:0] operation_194_2965;
reg [7:0] operation_194_2966_latch;
wire [7:0] operation_194_2966;
reg [7:0] operation_194_2967_latch;
wire [7:0] operation_194_2967;
reg [7:0] operation_194_2968_latch;
wire [7:0] operation_194_2968;
reg [7:0] operation_194_2969_latch;
wire [7:0] operation_194_2969;
reg [7:0] operation_194_2970_latch;
wire [7:0] operation_194_2970;
reg [7:0] operation_194_2971_latch;
wire [7:0] operation_194_2971;
reg [7:0] operation_194_2972_latch;
wire [7:0] operation_194_2972;
reg [7:0] operation_194_2973_latch;
wire [7:0] operation_194_2973;
reg [7:0] operation_194_2974_latch;
wire [7:0] operation_194_2974;
wire [7:0] operation_194_2128;
reg signed [31:0] operation_194_2129;
wire signed [31:0] operation_194_2130;
wire [7:0] operation_194_2132;
reg signed [31:0] operation_194_2133;
wire [7:0] operation_194_2134;
reg signed [31:0] operation_194_2135;
wire [7:0] operation_194_2136;
reg signed [31:0] operation_194_2137;
wire [7:0] operation_194_2138;
reg signed [31:0] operation_194_2139;
wire [7:0] operation_194_2140;
reg signed [31:0] operation_194_2141;
wire [7:0] operation_194_2142;
reg signed [31:0] operation_194_2143;
wire [7:0] operation_194_2144;
reg signed [31:0] operation_194_2145;
wire [7:0] operation_194_2146;
reg signed [31:0] operation_194_2147;
wire signed [31:0] operation_194_2148;
wire signed [31:0] operation_194_2149;
wire signed [31:0] operation_194_2150;
wire signed [31:0] operation_194_2151;
wire signed [31:0] operation_194_2152;
wire signed [31:0] operation_194_2153;
wire signed [31:0] operation_194_2154;
wire signed [31:0] operation_194_2155;
wire signed [31:0] operation_194_2156;
wire signed [31:0] operation_194_2157;
wire [7:0] operation_194_2158;
reg signed [31:0] operation_194_2159;
wire [7:0] operation_194_2160;
reg signed [31:0] operation_194_2161;
wire [7:0] operation_194_2162;
reg signed [31:0] operation_194_2163;
wire [7:0] operation_194_2164;
reg signed [31:0] operation_194_2165;
wire [7:0] operation_194_2166;
reg signed [31:0] operation_194_2167;
wire [7:0] operation_194_2168;
reg signed [31:0] operation_194_2169;
wire [7:0] operation_194_2170;
reg signed [31:0] operation_194_2171;
wire [7:0] operation_194_2172;
reg signed [31:0] operation_194_2173;
wire [7:0] operation_194_2174;
reg signed [31:0] operation_194_2175;
wire [7:0] operation_194_2176;
reg signed [31:0] operation_194_2177;
wire [7:0] operation_194_2178;
reg signed [31:0] operation_194_2179;
wire [7:0] operation_194_2180;
reg signed [31:0] operation_194_2181;
wire [7:0] operation_194_2182;
reg signed [31:0] operation_194_2183;
wire [7:0] operation_194_2184;
reg signed [31:0] operation_194_2185;
wire [7:0] operation_194_2186;
reg signed [31:0] operation_194_2187;
wire [7:0] operation_194_2188;
reg signed [31:0] operation_194_2189;
wire signed [31:0] operation_194_2190;
wire signed [31:0] operation_194_2191;
wire signed [31:0] operation_194_2192;
wire signed [31:0] operation_194_2193;
wire signed [31:0] operation_194_2194;
wire signed [31:0] operation_194_2195;
wire signed [31:0] operation_194_2196;
wire signed [31:0] operation_194_2197;
wire signed [31:0] operation_194_2198;
wire signed [31:0] operation_194_2199;
wire signed [31:0] operation_194_2200;
wire signed [31:0] operation_194_2201;
wire signed [31:0] operation_194_2202;
wire signed [31:0] operation_194_2203;
wire signed [31:0] operation_194_2204;
wire signed [31:0] operation_194_2205;
wire signed [31:0] operation_194_2206;
wire signed [31:0] operation_194_2207;
wire [7:0] operation_194_2208;
reg signed [31:0] operation_194_2209;
wire [7:0] operation_194_2210;
reg signed [31:0] operation_194_2211;
wire [7:0] operation_194_2212;
reg signed [31:0] operation_194_2213;
wire [7:0] operation_194_2214;
reg signed [31:0] operation_194_2215;
wire [7:0] operation_194_2216;
reg signed [31:0] operation_194_2217;
wire [7:0] operation_194_2218;
reg signed [31:0] operation_194_2219;
wire [7:0] operation_194_2220;
reg signed [31:0] operation_194_2221;
wire [7:0] operation_194_2222;
reg signed [31:0] operation_194_2223;
wire [7:0] operation_194_2224;
reg signed [31:0] operation_194_2225;
wire [7:0] operation_194_2226;
reg signed [31:0] operation_194_2227;
wire signed [31:0] operation_194_2228;
wire signed [31:0] operation_194_2229;
wire signed [31:0] operation_194_2230;
wire signed [31:0] operation_194_2231;
wire signed [31:0] operation_194_2232;
wire signed [31:0] operation_194_2233;
wire signed [31:0] operation_194_2234;
wire signed [31:0] operation_194_2235;
wire signed [31:0] operation_194_2236;
wire signed [31:0] operation_194_2237;
wire [7:0] operation_194_2238;
reg signed [31:0] operation_194_2239;
wire [7:0] operation_194_2240;
reg signed [31:0] operation_194_2241;
wire [7:0] operation_194_2242;
reg signed [31:0] operation_194_2243;
wire [7:0] operation_194_2244;
reg signed [31:0] operation_194_2245;
wire [7:0] operation_194_2246;
reg signed [31:0] operation_194_2247;
wire [7:0] operation_194_2248;
reg signed [31:0] operation_194_2249;
wire [7:0] operation_194_2250;
reg signed [31:0] operation_194_2251;
wire [7:0] operation_194_2252;
reg signed [31:0] operation_194_2253;
wire [7:0] operation_194_2254;
reg signed [31:0] operation_194_2255;
wire [7:0] operation_194_2256;
reg signed [31:0] operation_194_2257;
wire signed [31:0] operation_194_2258;
wire signed [31:0] operation_194_2259;
wire signed [31:0] operation_194_2260;
wire signed [31:0] operation_194_2261;
wire signed [31:0] operation_194_2262;
wire signed [31:0] operation_194_2263;
wire signed [31:0] operation_194_2264;
wire signed [31:0] operation_194_2265;
wire signed [31:0] operation_194_2266;
wire signed [31:0] operation_194_2267;
wire [7:0] operation_194_2268;
reg signed [31:0] operation_194_2269;
wire [7:0] operation_194_2270;
reg signed [31:0] operation_194_2271;
wire [7:0] operation_194_2272;
reg signed [31:0] operation_194_2273;
wire [7:0] operation_194_2274;
reg signed [31:0] operation_194_2275;
wire [7:0] operation_194_2276;
reg signed [31:0] operation_194_2277;
wire [7:0] operation_194_2278;
reg signed [31:0] operation_194_2279;
wire [7:0] operation_194_2280;
reg signed [31:0] operation_194_2281;
wire [7:0] operation_194_2282;
reg signed [31:0] operation_194_2283;
wire [7:0] operation_194_2284;
reg signed [31:0] operation_194_2285;
wire [7:0] operation_194_2286;
reg signed [31:0] operation_194_2287;
wire signed [31:0] operation_194_2288;
wire signed [31:0] operation_194_2289;
wire signed [31:0] operation_194_2290;
wire signed [31:0] operation_194_2291;
wire signed [31:0] operation_194_2292;
wire signed [31:0] operation_194_2293;
wire signed [31:0] operation_194_2294;
wire signed [31:0] operation_194_2295;
wire signed [31:0] operation_194_2296;
wire signed [31:0] operation_194_2297;
wire [7:0] operation_194_2298;
reg signed [31:0] operation_194_2299;
reg signed [31:0] operation_194_2300;
wire [7:0] operation_194_2301;
reg signed [31:0] operation_194_2302;
reg signed [31:0] operation_194_2303;
wire [7:0] operation_194_2304;
reg signed [31:0] operation_194_2305;
reg signed [31:0] operation_194_2306;
wire [7:0] operation_194_2307;
reg signed [31:0] operation_194_2308;
reg signed [31:0] operation_194_2309;
wire [7:0] operation_194_2310;
reg signed [31:0] operation_194_2311;
reg signed [31:0] operation_194_2312;
wire [7:0] operation_194_2313;
reg signed [31:0] operation_194_2314;
reg signed [31:0] operation_194_2315;
wire [7:0] operation_194_2316;
reg signed [31:0] operation_194_2317;
reg signed [31:0] operation_194_2318;
wire [7:0] operation_194_2319;
reg signed [31:0] operation_194_2320;
reg signed [31:0] operation_194_2321;
wire [7:0] operation_194_2322;
reg signed [31:0] operation_194_2323;
wire [7:0] operation_194_2324;
reg signed [31:0] operation_194_2325;
wire signed [31:0] operation_194_2326;
wire signed [31:0] operation_194_2327;
reg signed [31:0] operation_194_2328;
reg signed [31:0] operation_194_2329;
reg signed [31:0] operation_194_2330;
wire signed [31:0] operation_194_2331;
reg signed [31:0] operation_194_2332;
reg signed [31:0] operation_194_2333;
reg signed [31:0] operation_194_2334;
wire signed [31:0] operation_194_2335;
reg signed [31:0] operation_194_2336;
reg signed [31:0] operation_194_2337;
reg signed [31:0] operation_194_2338;
wire signed [31:0] operation_194_2339;
reg signed [31:0] operation_194_2340;
reg signed [31:0] operation_194_2341;
reg signed [31:0] operation_194_2342;
wire signed [31:0] operation_194_2343;
reg signed [31:0] operation_194_2344;
reg signed [31:0] operation_194_2345;
reg signed [31:0] operation_194_2346;
wire signed [31:0] operation_194_2347;
reg signed [31:0] operation_194_2348;
reg signed [31:0] operation_194_2349;
reg signed [31:0] operation_194_2350;
wire signed [31:0] operation_194_2351;
reg signed [31:0] operation_194_2352;
reg signed [31:0] operation_194_2353;
reg signed [31:0] operation_194_2354;
wire signed [31:0] operation_194_2355;
reg signed [31:0] operation_194_2356;
reg signed [31:0] operation_194_2357;
reg signed [31:0] operation_194_2358;
wire signed [31:0] operation_194_2359;
wire [7:0] operation_194_2360;
reg signed [31:0] operation_194_2361;
reg signed [31:0] operation_194_2362;
wire [7:0] operation_194_2363;
reg signed [31:0] operation_194_2364;
reg signed [31:0] operation_194_2365;
wire [7:0] operation_194_2366;
reg signed [31:0] operation_194_2367;
reg signed [31:0] operation_194_2368;
wire [7:0] operation_194_2369;
reg signed [31:0] operation_194_2370;
reg signed [31:0] operation_194_2371;
wire [7:0] operation_194_2372;
reg signed [31:0] operation_194_2373;
reg signed [31:0] operation_194_2374;
wire [7:0] operation_194_2375;
reg signed [31:0] operation_194_2376;
reg signed [31:0] operation_194_2377;
wire [7:0] operation_194_2378;
reg signed [31:0] operation_194_2379;
reg signed [31:0] operation_194_2380;
wire [7:0] operation_194_2381;
reg signed [31:0] operation_194_2382;
reg signed [31:0] operation_194_2383;
wire [7:0] operation_194_2384;
reg signed [31:0] operation_194_2385;
wire [7:0] operation_194_2386;
reg signed [31:0] operation_194_2387;
wire signed [31:0] operation_194_2388;
wire signed [31:0] operation_194_2389;
wire signed [31:0] operation_194_2390;
wire signed [31:0] operation_194_2391;
reg signed [31:0] operation_194_2392;
reg signed [31:0] operation_194_2393;
reg signed [31:0] operation_194_2394;
wire signed [31:0] operation_194_2395;
reg signed [31:0] operation_194_2396;
reg signed [31:0] operation_194_2397;
reg signed [31:0] operation_194_2398;
wire signed [31:0] operation_194_2399;
reg signed [31:0] operation_194_2400;
reg signed [31:0] operation_194_2401;
reg signed [31:0] operation_194_2402;
wire signed [31:0] operation_194_2403;
reg signed [31:0] operation_194_2404;
reg signed [31:0] operation_194_2405;
reg signed [31:0] operation_194_2406;
wire signed [31:0] operation_194_2407;
reg signed [31:0] operation_194_2408;
reg signed [31:0] operation_194_2409;
reg signed [31:0] operation_194_2410;
wire signed [31:0] operation_194_2411;
reg signed [31:0] operation_194_2412;
reg signed [31:0] operation_194_2413;
reg signed [31:0] operation_194_2414;
wire signed [31:0] operation_194_2415;
reg signed [31:0] operation_194_2416;
reg signed [31:0] operation_194_2417;
reg signed [31:0] operation_194_2418;
wire signed [31:0] operation_194_2419;
reg signed [31:0] operation_194_2420;
reg signed [31:0] operation_194_2421;
reg signed [31:0] operation_194_2422;
wire signed [31:0] operation_194_2423;
wire [7:0] operation_194_2424;
wire [7:0] operation_194_2425;
reg signed [31:0] operation_194_2426;
wire [7:0] operation_194_2427;
wire [7:0] operation_194_2428;
reg signed [31:0] operation_194_2429;
wire [7:0] operation_194_2430;
wire [7:0] operation_194_2431;
reg signed [31:0] operation_194_2432;
wire [7:0] operation_194_2433;
wire [7:0] operation_194_2434;
reg signed [31:0] operation_194_2435;
wire [7:0] operation_194_2436;
reg signed [31:0] operation_194_2437;
wire [7:0] operation_194_2438;
reg signed [31:0] operation_194_2439;
wire [7:0] operation_194_2440;
reg signed [31:0] operation_194_2441;
wire [7:0] operation_194_2442;
reg signed [31:0] operation_194_2443;
wire [7:0] operation_194_2444;
reg signed [31:0] operation_194_2445;
wire signed [31:0] operation_194_2446;
wire signed [31:0] operation_194_2447;
wire signed [31:0] operation_194_2448;
wire signed [31:0] operation_194_2449;
wire signed [31:0] operation_194_2450;
reg signed [31:0] operation_194_2451;
reg signed [31:0] operation_194_2452;
reg signed [31:0] operation_194_2453;
reg signed [31:0] operation_194_2454;
wire [7:0] operation_194_2455;
reg signed [31:0] operation_194_2456;
wire [7:0] operation_194_2457;
reg signed [31:0] operation_194_2458;
wire [7:0] operation_194_2459;
reg signed [31:0] operation_194_2460;
wire [7:0] operation_194_2461;
reg signed [31:0] operation_194_2462;
wire [7:0] operation_194_2463;
reg signed [31:0] operation_194_2464;
wire [7:0] operation_194_2465;
reg signed [31:0] operation_194_2466;
wire [7:0] operation_194_2467;
reg signed [31:0] operation_194_2468;
wire [7:0] operation_194_2469;
reg signed [31:0] operation_194_2470;
wire [7:0] operation_194_2471;
reg signed [31:0] operation_194_2472;
wire [7:0] operation_194_2473;
reg signed [31:0] operation_194_2474;
wire [7:0] operation_194_2475;
reg signed [31:0] operation_194_2476;
wire signed [31:0] operation_194_2483;
reg signed [31:0] operation_194_2486;
reg signed [31:0] operation_194_2487;
reg signed [31:0] operation_194_2488;
reg signed [31:0] operation_194_2489;
wire signed [31:0] operation_194_2490;
wire signed [31:0] operation_194_2491;
wire signed [31:0] operation_194_2492;
wire signed [31:0] operation_194_2493;
wire signed [31:0] operation_194_2494;
wire signed [31:0] operation_194_2495;
wire signed [31:0] operation_194_2496;
wire signed [31:0] operation_194_2497;
wire [7:0] operation_194_2500;
reg signed [31:0] operation_194_2501;
wire [7:0] operation_194_2502;
reg signed [31:0] operation_194_2503;
wire signed [31:0] operation_194_2514;
wire signed [31:0] operation_194_2516;
reg [7:0] operation_194_2518_latch;
wire [7:0] operation_194_2518;
reg [7:0] operation_194_2519_latch;
wire [7:0] operation_194_2519;
wire signed [31:0] operation_194_2520;
wire signed [31:0] operation_194_2521;
wire signed [31:0] operation_194_2522;
wire signed [31:0] operation_194_2523;
wire signed [31:0] operation_194_2524;
wire signed [31:0] operation_194_2525;
wire signed [31:0] operation_194_2526;
wire signed [31:0] operation_194_2527;
reg [7:0] operation_194_2528_latch;
wire [7:0] operation_194_2528;
reg [7:0] operation_194_2529_latch;
wire [7:0] operation_194_2529;
reg [7:0] operation_194_2530_latch;
wire [7:0] operation_194_2530;
reg [7:0] operation_194_2531_latch;
wire [7:0] operation_194_2531;
reg [7:0] operation_194_2532_latch;
wire [7:0] operation_194_2532;
reg [7:0] operation_194_2533_latch;
wire [7:0] operation_194_2533;
reg [7:0] operation_194_2534_latch;
wire [7:0] operation_194_2534;
reg [7:0] operation_194_2535_latch;
wire [7:0] operation_194_2535;
reg [7:0] operation_194_2536_latch;
wire [7:0] operation_194_2536;
reg [7:0] operation_194_2537_latch;
wire [7:0] operation_194_2537;
reg [7:0] operation_194_2538_latch;
wire [7:0] operation_194_2538;
reg [7:0] operation_194_2539_latch;
wire [7:0] operation_194_2539;
reg [7:0] operation_194_2540_latch;
wire [7:0] operation_194_2540;
reg [7:0] operation_194_2541_latch;
wire [7:0] operation_194_2541;
reg [7:0] operation_194_2542_latch;
wire [7:0] operation_194_2542;
reg [7:0] operation_194_2543_latch;
wire [7:0] operation_194_2543;
reg [7:0] operation_194_2544_latch;
wire [7:0] operation_194_2544;
reg [7:0] operation_194_2545_latch;
wire [7:0] operation_194_2545;
wire [7:0] operation_194_1699;
reg signed [31:0] operation_194_1700;
wire signed [31:0] operation_194_1701;
wire [7:0] operation_194_1703;
reg signed [31:0] operation_194_1704;
wire [7:0] operation_194_1705;
reg signed [31:0] operation_194_1706;
wire [7:0] operation_194_1707;
reg signed [31:0] operation_194_1708;
wire [7:0] operation_194_1709;
reg signed [31:0] operation_194_1710;
wire [7:0] operation_194_1711;
reg signed [31:0] operation_194_1712;
wire [7:0] operation_194_1713;
reg signed [31:0] operation_194_1714;
wire [7:0] operation_194_1715;
reg signed [31:0] operation_194_1716;
wire [7:0] operation_194_1717;
reg signed [31:0] operation_194_1718;
wire signed [31:0] operation_194_1719;
wire signed [31:0] operation_194_1720;
wire signed [31:0] operation_194_1721;
wire signed [31:0] operation_194_1722;
wire signed [31:0] operation_194_1723;
wire signed [31:0] operation_194_1724;
wire signed [31:0] operation_194_1725;
wire signed [31:0] operation_194_1726;
wire signed [31:0] operation_194_1727;
wire signed [31:0] operation_194_1728;
wire [7:0] operation_194_1729;
reg signed [31:0] operation_194_1730;
wire [7:0] operation_194_1731;
reg signed [31:0] operation_194_1732;
wire [7:0] operation_194_1733;
reg signed [31:0] operation_194_1734;
wire [7:0] operation_194_1735;
reg signed [31:0] operation_194_1736;
wire [7:0] operation_194_1737;
reg signed [31:0] operation_194_1738;
wire [7:0] operation_194_1739;
reg signed [31:0] operation_194_1740;
wire [7:0] operation_194_1741;
reg signed [31:0] operation_194_1742;
wire [7:0] operation_194_1743;
reg signed [31:0] operation_194_1744;
wire [7:0] operation_194_1745;
reg signed [31:0] operation_194_1746;
wire [7:0] operation_194_1747;
reg signed [31:0] operation_194_1748;
wire [7:0] operation_194_1749;
reg signed [31:0] operation_194_1750;
wire [7:0] operation_194_1751;
reg signed [31:0] operation_194_1752;
wire [7:0] operation_194_1753;
reg signed [31:0] operation_194_1754;
wire [7:0] operation_194_1755;
reg signed [31:0] operation_194_1756;
wire [7:0] operation_194_1757;
reg signed [31:0] operation_194_1758;
wire [7:0] operation_194_1759;
reg signed [31:0] operation_194_1760;
wire signed [31:0] operation_194_1761;
wire signed [31:0] operation_194_1762;
wire signed [31:0] operation_194_1763;
wire signed [31:0] operation_194_1764;
wire signed [31:0] operation_194_1765;
wire signed [31:0] operation_194_1766;
wire signed [31:0] operation_194_1767;
wire signed [31:0] operation_194_1768;
wire signed [31:0] operation_194_1769;
wire signed [31:0] operation_194_1770;
wire signed [31:0] operation_194_1771;
wire signed [31:0] operation_194_1772;
wire signed [31:0] operation_194_1773;
wire signed [31:0] operation_194_1774;
wire signed [31:0] operation_194_1775;
wire signed [31:0] operation_194_1776;
wire signed [31:0] operation_194_1777;
wire signed [31:0] operation_194_1778;
wire [7:0] operation_194_1779;
reg signed [31:0] operation_194_1780;
wire [7:0] operation_194_1781;
reg signed [31:0] operation_194_1782;
wire [7:0] operation_194_1783;
reg signed [31:0] operation_194_1784;
wire [7:0] operation_194_1785;
reg signed [31:0] operation_194_1786;
wire [7:0] operation_194_1787;
reg signed [31:0] operation_194_1788;
wire [7:0] operation_194_1789;
reg signed [31:0] operation_194_1790;
wire [7:0] operation_194_1791;
reg signed [31:0] operation_194_1792;
wire [7:0] operation_194_1793;
reg signed [31:0] operation_194_1794;
wire [7:0] operation_194_1795;
reg signed [31:0] operation_194_1796;
wire [7:0] operation_194_1797;
reg signed [31:0] operation_194_1798;
wire signed [31:0] operation_194_1799;
wire signed [31:0] operation_194_1800;
wire signed [31:0] operation_194_1801;
wire signed [31:0] operation_194_1802;
wire signed [31:0] operation_194_1803;
wire signed [31:0] operation_194_1804;
wire signed [31:0] operation_194_1805;
wire signed [31:0] operation_194_1806;
wire signed [31:0] operation_194_1807;
wire signed [31:0] operation_194_1808;
wire [7:0] operation_194_1809;
reg signed [31:0] operation_194_1810;
wire [7:0] operation_194_1811;
reg signed [31:0] operation_194_1812;
wire [7:0] operation_194_1813;
reg signed [31:0] operation_194_1814;
wire [7:0] operation_194_1815;
reg signed [31:0] operation_194_1816;
wire [7:0] operation_194_1817;
reg signed [31:0] operation_194_1818;
wire [7:0] operation_194_1819;
reg signed [31:0] operation_194_1820;
wire [7:0] operation_194_1821;
reg signed [31:0] operation_194_1822;
wire [7:0] operation_194_1823;
reg signed [31:0] operation_194_1824;
wire [7:0] operation_194_1825;
reg signed [31:0] operation_194_1826;
wire [7:0] operation_194_1827;
reg signed [31:0] operation_194_1828;
wire signed [31:0] operation_194_1829;
wire signed [31:0] operation_194_1830;
wire signed [31:0] operation_194_1831;
wire signed [31:0] operation_194_1832;
wire signed [31:0] operation_194_1833;
wire signed [31:0] operation_194_1834;
wire signed [31:0] operation_194_1835;
wire signed [31:0] operation_194_1836;
wire signed [31:0] operation_194_1837;
wire signed [31:0] operation_194_1838;
wire [7:0] operation_194_1839;
reg signed [31:0] operation_194_1840;
wire [7:0] operation_194_1841;
reg signed [31:0] operation_194_1842;
wire [7:0] operation_194_1843;
reg signed [31:0] operation_194_1844;
wire [7:0] operation_194_1845;
reg signed [31:0] operation_194_1846;
wire [7:0] operation_194_1847;
reg signed [31:0] operation_194_1848;
wire [7:0] operation_194_1849;
reg signed [31:0] operation_194_1850;
wire [7:0] operation_194_1851;
reg signed [31:0] operation_194_1852;
wire [7:0] operation_194_1853;
reg signed [31:0] operation_194_1854;
wire [7:0] operation_194_1855;
reg signed [31:0] operation_194_1856;
wire [7:0] operation_194_1857;
reg signed [31:0] operation_194_1858;
wire signed [31:0] operation_194_1859;
wire signed [31:0] operation_194_1860;
wire signed [31:0] operation_194_1861;
wire signed [31:0] operation_194_1862;
wire signed [31:0] operation_194_1863;
wire signed [31:0] operation_194_1864;
wire signed [31:0] operation_194_1865;
wire signed [31:0] operation_194_1866;
wire signed [31:0] operation_194_1867;
wire signed [31:0] operation_194_1868;
wire [7:0] operation_194_1869;
reg signed [31:0] operation_194_1870;
reg signed [31:0] operation_194_1871;
wire [7:0] operation_194_1872;
reg signed [31:0] operation_194_1873;
reg signed [31:0] operation_194_1874;
wire [7:0] operation_194_1875;
reg signed [31:0] operation_194_1876;
reg signed [31:0] operation_194_1877;
wire [7:0] operation_194_1878;
reg signed [31:0] operation_194_1879;
reg signed [31:0] operation_194_1880;
wire [7:0] operation_194_1881;
reg signed [31:0] operation_194_1882;
reg signed [31:0] operation_194_1883;
wire [7:0] operation_194_1884;
reg signed [31:0] operation_194_1885;
reg signed [31:0] operation_194_1886;
wire [7:0] operation_194_1887;
reg signed [31:0] operation_194_1888;
reg signed [31:0] operation_194_1889;
wire [7:0] operation_194_1890;
reg signed [31:0] operation_194_1891;
reg signed [31:0] operation_194_1892;
wire [7:0] operation_194_1893;
reg signed [31:0] operation_194_1894;
wire [7:0] operation_194_1895;
reg signed [31:0] operation_194_1896;
wire signed [31:0] operation_194_1897;
wire signed [31:0] operation_194_1898;
reg signed [31:0] operation_194_1899;
reg signed [31:0] operation_194_1900;
reg signed [31:0] operation_194_1901;
wire signed [31:0] operation_194_1902;
reg signed [31:0] operation_194_1903;
reg signed [31:0] operation_194_1904;
reg signed [31:0] operation_194_1905;
wire signed [31:0] operation_194_1906;
reg signed [31:0] operation_194_1907;
reg signed [31:0] operation_194_1908;
reg signed [31:0] operation_194_1909;
wire signed [31:0] operation_194_1910;
reg signed [31:0] operation_194_1911;
reg signed [31:0] operation_194_1912;
reg signed [31:0] operation_194_1913;
wire signed [31:0] operation_194_1914;
reg signed [31:0] operation_194_1915;
reg signed [31:0] operation_194_1916;
reg signed [31:0] operation_194_1917;
wire signed [31:0] operation_194_1918;
reg signed [31:0] operation_194_1919;
reg signed [31:0] operation_194_1920;
reg signed [31:0] operation_194_1921;
wire signed [31:0] operation_194_1922;
reg signed [31:0] operation_194_1923;
reg signed [31:0] operation_194_1924;
reg signed [31:0] operation_194_1925;
wire signed [31:0] operation_194_1926;
reg signed [31:0] operation_194_1927;
reg signed [31:0] operation_194_1928;
reg signed [31:0] operation_194_1929;
wire signed [31:0] operation_194_1930;
wire [7:0] operation_194_1931;
reg signed [31:0] operation_194_1932;
reg signed [31:0] operation_194_1933;
wire [7:0] operation_194_1934;
reg signed [31:0] operation_194_1935;
reg signed [31:0] operation_194_1936;
wire [7:0] operation_194_1937;
reg signed [31:0] operation_194_1938;
reg signed [31:0] operation_194_1939;
wire [7:0] operation_194_1940;
reg signed [31:0] operation_194_1941;
reg signed [31:0] operation_194_1942;
wire [7:0] operation_194_1943;
reg signed [31:0] operation_194_1944;
reg signed [31:0] operation_194_1945;
wire [7:0] operation_194_1946;
reg signed [31:0] operation_194_1947;
reg signed [31:0] operation_194_1948;
wire [7:0] operation_194_1949;
reg signed [31:0] operation_194_1950;
reg signed [31:0] operation_194_1951;
wire [7:0] operation_194_1952;
reg signed [31:0] operation_194_1953;
reg signed [31:0] operation_194_1954;
wire [7:0] operation_194_1955;
reg signed [31:0] operation_194_1956;
wire [7:0] operation_194_1957;
reg signed [31:0] operation_194_1958;
wire signed [31:0] operation_194_1959;
wire signed [31:0] operation_194_1960;
wire signed [31:0] operation_194_1961;
wire signed [31:0] operation_194_1962;
reg signed [31:0] operation_194_1963;
reg signed [31:0] operation_194_1964;
reg signed [31:0] operation_194_1965;
wire signed [31:0] operation_194_1966;
reg signed [31:0] operation_194_1967;
reg signed [31:0] operation_194_1968;
reg signed [31:0] operation_194_1969;
wire signed [31:0] operation_194_1970;
reg signed [31:0] operation_194_1971;
reg signed [31:0] operation_194_1972;
reg signed [31:0] operation_194_1973;
wire signed [31:0] operation_194_1974;
reg signed [31:0] operation_194_1975;
reg signed [31:0] operation_194_1976;
reg signed [31:0] operation_194_1977;
wire signed [31:0] operation_194_1978;
reg signed [31:0] operation_194_1979;
reg signed [31:0] operation_194_1980;
reg signed [31:0] operation_194_1981;
wire signed [31:0] operation_194_1982;
reg signed [31:0] operation_194_1983;
reg signed [31:0] operation_194_1984;
reg signed [31:0] operation_194_1985;
wire signed [31:0] operation_194_1986;
reg signed [31:0] operation_194_1987;
reg signed [31:0] operation_194_1988;
reg signed [31:0] operation_194_1989;
wire signed [31:0] operation_194_1990;
reg signed [31:0] operation_194_1991;
reg signed [31:0] operation_194_1992;
reg signed [31:0] operation_194_1993;
wire signed [31:0] operation_194_1994;
wire [7:0] operation_194_1995;
wire [7:0] operation_194_1996;
reg signed [31:0] operation_194_1997;
wire [7:0] operation_194_1998;
wire [7:0] operation_194_1999;
reg signed [31:0] operation_194_2000;
wire [7:0] operation_194_2001;
wire [7:0] operation_194_2002;
reg signed [31:0] operation_194_2003;
wire [7:0] operation_194_2004;
wire [7:0] operation_194_2005;
reg signed [31:0] operation_194_2006;
wire [7:0] operation_194_2007;
reg signed [31:0] operation_194_2008;
wire [7:0] operation_194_2009;
reg signed [31:0] operation_194_2010;
wire [7:0] operation_194_2011;
reg signed [31:0] operation_194_2012;
wire [7:0] operation_194_2013;
reg signed [31:0] operation_194_2014;
wire [7:0] operation_194_2015;
reg signed [31:0] operation_194_2016;
wire signed [31:0] operation_194_2017;
wire signed [31:0] operation_194_2018;
wire signed [31:0] operation_194_2019;
wire signed [31:0] operation_194_2020;
wire signed [31:0] operation_194_2021;
reg signed [31:0] operation_194_2022;
reg signed [31:0] operation_194_2023;
reg signed [31:0] operation_194_2024;
reg signed [31:0] operation_194_2025;
wire [7:0] operation_194_2026;
reg signed [31:0] operation_194_2027;
wire [7:0] operation_194_2028;
reg signed [31:0] operation_194_2029;
wire [7:0] operation_194_2030;
reg signed [31:0] operation_194_2031;
wire [7:0] operation_194_2032;
reg signed [31:0] operation_194_2033;
wire [7:0] operation_194_2034;
reg signed [31:0] operation_194_2035;
wire [7:0] operation_194_2036;
reg signed [31:0] operation_194_2037;
wire [7:0] operation_194_2038;
reg signed [31:0] operation_194_2039;
wire [7:0] operation_194_2040;
reg signed [31:0] operation_194_2041;
wire [7:0] operation_194_2042;
reg signed [31:0] operation_194_2043;
wire [7:0] operation_194_2044;
reg signed [31:0] operation_194_2045;
wire [7:0] operation_194_2046;
reg signed [31:0] operation_194_2047;
wire signed [31:0] operation_194_2054;
reg signed [31:0] operation_194_2057;
reg signed [31:0] operation_194_2058;
reg signed [31:0] operation_194_2059;
reg signed [31:0] operation_194_2060;
wire signed [31:0] operation_194_2061;
wire signed [31:0] operation_194_2062;
wire signed [31:0] operation_194_2063;
wire signed [31:0] operation_194_2064;
wire signed [31:0] operation_194_2065;
wire signed [31:0] operation_194_2066;
wire signed [31:0] operation_194_2067;
wire signed [31:0] operation_194_2068;
wire [7:0] operation_194_2071;
reg signed [31:0] operation_194_2072;
wire [7:0] operation_194_2073;
reg signed [31:0] operation_194_2074;
wire signed [31:0] operation_194_2085;
wire signed [31:0] operation_194_2087;
reg [7:0] operation_194_2089_latch;
wire [7:0] operation_194_2089;
reg [7:0] operation_194_2090_latch;
wire [7:0] operation_194_2090;
wire signed [31:0] operation_194_2091;
wire signed [31:0] operation_194_2092;
wire signed [31:0] operation_194_2093;
wire signed [31:0] operation_194_2094;
wire signed [31:0] operation_194_2095;
wire signed [31:0] operation_194_2096;
wire signed [31:0] operation_194_2097;
wire signed [31:0] operation_194_2098;
reg [7:0] operation_194_2099_latch;
wire [7:0] operation_194_2099;
reg [7:0] operation_194_2100_latch;
wire [7:0] operation_194_2100;
reg [7:0] operation_194_2101_latch;
wire [7:0] operation_194_2101;
reg [7:0] operation_194_2102_latch;
wire [7:0] operation_194_2102;
reg [7:0] operation_194_2103_latch;
wire [7:0] operation_194_2103;
reg [7:0] operation_194_2104_latch;
wire [7:0] operation_194_2104;
reg [7:0] operation_194_2105_latch;
wire [7:0] operation_194_2105;
reg [7:0] operation_194_2106_latch;
wire [7:0] operation_194_2106;
reg [7:0] operation_194_2107_latch;
wire [7:0] operation_194_2107;
reg [7:0] operation_194_2108_latch;
wire [7:0] operation_194_2108;
reg [7:0] operation_194_2109_latch;
wire [7:0] operation_194_2109;
reg [7:0] operation_194_2110_latch;
wire [7:0] operation_194_2110;
reg [7:0] operation_194_2111_latch;
wire [7:0] operation_194_2111;
reg [7:0] operation_194_2112_latch;
wire [7:0] operation_194_2112;
reg [7:0] operation_194_2113_latch;
wire [7:0] operation_194_2113;
reg [7:0] operation_194_2114_latch;
wire [7:0] operation_194_2114;
reg [7:0] operation_194_2115_latch;
wire [7:0] operation_194_2115;
reg [7:0] operation_194_2116_latch;
wire [7:0] operation_194_2116;
wire [7:0] operation_194_127;
reg signed [31:0] operation_194_126;
wire signed [31:0] operation_194_123;
wire [7:0] operation_194_7;
reg signed [31:0] operation_194_6;
wire [7:0] operation_194_23;
reg signed [31:0] operation_194_22;
wire [7:0] operation_194_39;
reg signed [31:0] operation_194_38;
wire [7:0] operation_194_55;
reg signed [31:0] operation_194_54;
wire [7:0] operation_194_71;
reg signed [31:0] operation_194_70;
wire [7:0] operation_194_87;
reg signed [31:0] operation_194_86;
wire [7:0] operation_194_103;
reg signed [31:0] operation_194_102;
wire [7:0] operation_194_119;
reg signed [31:0] operation_194_118;
wire signed [31:0] operation_194_117;
wire signed [31:0] operation_194_115;
wire signed [31:0] operation_194_101;
wire signed [31:0] operation_194_99;
wire signed [31:0] operation_194_85;
wire signed [31:0] operation_194_83;
wire signed [31:0] operation_194_69;
wire signed [31:0] operation_194_67;
wire signed [31:0] operation_194_53;
wire signed [31:0] operation_194_51;
wire signed [31:0] operation_194_37;
wire signed [31:0] operation_194_35;
wire signed [31:0] operation_194_21;
wire signed [31:0] operation_194_19;
wire signed [31:0] operation_194_5;
wire signed [31:0] operation_194_3;
wire [7:0] operation_194_15;
reg signed [31:0] operation_194_14;
wire signed [31:0] operation_194_11;
wire signed [31:0] operation_194_13;
wire [7:0] operation_194_31;
reg signed [31:0] operation_194_30;
wire signed [31:0] operation_194_27;
wire signed [31:0] operation_194_29;
wire [7:0] operation_194_47;
reg signed [31:0] operation_194_46;
wire signed [31:0] operation_194_43;
wire signed [31:0] operation_194_45;
wire [7:0] operation_194_63;
reg signed [31:0] operation_194_62;
wire signed [31:0] operation_194_59;
wire signed [31:0] operation_194_61;
wire [7:0] operation_194_79;
reg signed [31:0] operation_194_78;
wire signed [31:0] operation_194_75;
wire signed [31:0] operation_194_77;
wire [7:0] operation_194_95;
reg signed [31:0] operation_194_94;
wire signed [31:0] operation_194_91;
wire signed [31:0] operation_194_93;
wire [7:0] operation_194_111;
reg signed [31:0] operation_194_110;
wire signed [31:0] operation_194_107;
wire signed [31:0] operation_194_109;
wire signed [31:0] operation_194_125;
wire signed [31:0] operation_194_5601;
wire signed [31:0] operation_194_5597;
wire signed [31:0] operation_194_5592;
wire signed [31:0] operation_194_5587;
wire signed [31:0] operation_194_5582;
wire signed [31:0] operation_194_5577;
wire signed [31:0] operation_194_5572;
wire signed [31:0] operation_194_5567;
wire signed [31:0] operation_194_5562;
wire signed [31:0] operation_194_5557;
wire signed [31:0] operation_194_2119;
wire [127:0] operation_194_124;
wire [127:0] operation_194_122;
reg control_194_follow;
wire control_194_end;
wire control_194_0;
reg control_194_start;
reg control_194_83;
reg control_194_82;
reg control_194_81;
reg control_194_80;
reg control_194_79;
reg control_194_78;
reg control_194_77;
reg control_194_76;
reg control_194_75;
reg control_194_74;
reg control_194_73;
reg control_194_72;
reg control_194_71;
reg control_194_70;
reg control_194_69;
reg control_194_68;
reg control_194_67;
reg control_194_66;
reg control_194_65;
reg control_194_64;
reg control_194_63;
reg control_194_62;
reg control_194_61;
reg control_194_60;
reg control_194_59;
reg control_194_58;
reg control_194_57;
reg control_194_56;
reg control_194_55;
reg control_194_54;
reg control_194_53;
reg control_194_52;
reg control_194_51;
reg control_194_50;
reg control_194_49;
reg control_194_48;
reg control_194_47;
reg control_194_46;
reg control_194_45;
reg control_194_44;
reg control_194_43;
reg control_194_42;
reg control_194_41;
reg control_194_40;
reg control_194_39;
reg control_194_38;
reg control_194_37;
reg control_194_36;
reg control_194_35;
reg control_194_34;
reg control_194_33;
reg control_194_32;
reg control_194_31;
reg control_194_30;
reg control_194_29;
reg control_194_28;
reg control_194_27;
reg control_194_26;
reg control_194_25;
reg control_194_24;
reg control_194_23;
reg control_194_22;
reg control_194_21;
reg control_194_20;
reg control_194_19;
reg control_194_18;
reg control_194_17;
reg control_194_16;
reg control_194_15;
reg control_194_14;
reg control_194_13;
reg control_194_12;
reg control_194_11;
reg control_194_10;
reg control_194_9;
reg control_194_8;
reg control_194_7;
reg control_194_6;
reg control_194_5;
reg control_194_4;
reg control_194_3;
reg control_194_2;
reg control_194_1;
reg [127:0] input_key_194_follow;
wire [127:0] input_key_194;
reg [127:0] input_in_194_follow;
wire [127:0] input_in_194;
reg [7:0] lookup_sbox_0_output;
reg [7:0] sbox_0[256];
wire lookup_sbox_0_enable;
wire [255:0] lookup_sbox_0_0;
reg [7:0] lookup_sbox_1_output;
reg [7:0] sbox_1[256];
wire lookup_sbox_1_enable;
wire [255:0] lookup_sbox_1_0;
reg [7:0] lookup_sbox_2_output;
reg [7:0] sbox_2[256];
wire lookup_sbox_2_enable;
wire [255:0] lookup_sbox_2_0;
reg [7:0] lookup_sbox_3_output;
reg [7:0] sbox_3[256];
wire lookup_sbox_3_enable;
wire [255:0] lookup_sbox_3_0;
reg [7:0] lookup_sbox_4_output;
reg [7:0] sbox_4[256];
wire lookup_sbox_4_enable;
wire [255:0] lookup_sbox_4_0;
reg [7:0] lookup_sbox_5_output;
reg [7:0] sbox_5[256];
wire lookup_sbox_5_enable;
wire [255:0] lookup_sbox_5_0;
reg [7:0] lookup_sbox_6_output;
reg [7:0] sbox_6[256];
wire lookup_sbox_6_enable;
wire [255:0] lookup_sbox_6_0;
reg [7:0] lookup_sbox_7_output;
reg [7:0] sbox_7[256];
wire lookup_sbox_7_enable;
wire [255:0] lookup_sbox_7_0;
reg [7:0] lookup_sbox_8_output;
reg [7:0] sbox_8[256];
wire lookup_sbox_8_enable;
wire [255:0] lookup_sbox_8_0;
reg [7:0] lookup_sbox_9_output;
reg [7:0] sbox_9[256];
wire lookup_sbox_9_enable;
wire [255:0] lookup_sbox_9_0;
reg [7:0] lookup_sbox_10_output;
reg [7:0] sbox_10[256];
wire lookup_sbox_10_enable;
wire [255:0] lookup_sbox_10_0;
reg [7:0] lookup_sbox_11_output;
reg [7:0] sbox_11[256];
wire lookup_sbox_11_enable;
wire [255:0] lookup_sbox_11_0;
reg [7:0] lookup_sbox_12_output;
reg [7:0] sbox_12[256];
wire lookup_sbox_12_enable;
wire [255:0] lookup_sbox_12_0;
reg [7:0] lookup_sbox_13_output;
reg [7:0] sbox_13[256];
wire lookup_sbox_13_enable;
wire [255:0] lookup_sbox_13_0;
reg [7:0] lookup_sbox_14_output;
reg [7:0] sbox_14[256];
wire lookup_sbox_14_enable;
wire [255:0] lookup_sbox_14_0;
reg [7:0] lookup_sbox_15_output;
reg [7:0] sbox_15[256];
wire lookup_sbox_15_enable;
wire [255:0] lookup_sbox_15_0;
reg [7:0] lookup_sbox_16_output;
reg [7:0] sbox_16[256];
wire lookup_sbox_16_enable;
wire [255:0] lookup_sbox_16_0;
reg [7:0] lookup_sbox_17_output;
reg [7:0] sbox_17[256];
wire lookup_sbox_17_enable;
wire [255:0] lookup_sbox_17_0;
reg [7:0] lookup_sbox_18_output;
reg [7:0] sbox_18[256];
wire lookup_sbox_18_enable;
wire [255:0] lookup_sbox_18_0;
reg [7:0] lookup_sbox_19_output;
reg [7:0] sbox_19[256];
wire lookup_sbox_19_enable;
wire [255:0] lookup_sbox_19_0;
reg [7:0] lookup_sbox_20_output;
reg [7:0] sbox_20[256];
wire lookup_sbox_20_enable;
wire [255:0] lookup_sbox_20_0;
reg [7:0] lookup_sbox_21_output;
reg [7:0] sbox_21[256];
wire lookup_sbox_21_enable;
wire [255:0] lookup_sbox_21_0;
reg [7:0] lookup_sbox_22_output;
reg [7:0] sbox_22[256];
wire lookup_sbox_22_enable;
wire [255:0] lookup_sbox_22_0;
reg [7:0] lookup_sbox_23_output;
reg [7:0] sbox_23[256];
wire lookup_sbox_23_enable;
wire [255:0] lookup_sbox_23_0;
reg [7:0] lookup_sbox_24_output;
reg [7:0] sbox_24[256];
wire lookup_sbox_24_enable;
wire [255:0] lookup_sbox_24_0;
reg [7:0] lookup_sbox_25_output;
reg [7:0] sbox_25[256];
wire lookup_sbox_25_enable;
wire [255:0] lookup_sbox_25_0;
reg [7:0] lookup_sbox_26_output;
reg [7:0] sbox_26[256];
wire lookup_sbox_26_enable;
wire [255:0] lookup_sbox_26_0;
reg [7:0] lookup_sbox_27_output;
reg [7:0] sbox_27[256];
wire lookup_sbox_27_enable;
wire [255:0] lookup_sbox_27_0;
reg [7:0] lookup_sbox_28_output;
reg [7:0] sbox_28[256];
wire lookup_sbox_28_enable;
wire [255:0] lookup_sbox_28_0;
reg [7:0] lookup_sbox_29_output;
reg [7:0] sbox_29[256];
wire lookup_sbox_29_enable;
wire [255:0] lookup_sbox_29_0;
reg [7:0] lookup_sbox_30_output;
reg [7:0] sbox_30[256];
wire lookup_sbox_30_enable;
wire [255:0] lookup_sbox_30_0;
reg [7:0] lookup_sbox_31_output;
reg [7:0] sbox_31[256];
wire lookup_sbox_31_enable;
wire [255:0] lookup_sbox_31_0;
reg startfollow;
initial begin
    
    sbox_0[0] = 8'd99;
    sbox_0[1] = 8'd124;
    sbox_0[2] = 8'd119;
    sbox_0[3] = 8'd123;
    sbox_0[4] = 8'd242;
    sbox_0[5] = 8'd107;
    sbox_0[6] = 8'd111;
    sbox_0[7] = 8'd197;
    sbox_0[8] = 8'd48;
    sbox_0[9] = 8'd1;
    sbox_0[10] = 8'd103;
    sbox_0[11] = 8'd43;
    sbox_0[12] = 8'd254;
    sbox_0[13] = 8'd215;
    sbox_0[14] = 8'd171;
    sbox_0[15] = 8'd118;
    sbox_0[16] = 8'd202;
    sbox_0[17] = 8'd130;
    sbox_0[18] = 8'd201;
    sbox_0[19] = 8'd125;
    sbox_0[20] = 8'd250;
    sbox_0[21] = 8'd89;
    sbox_0[22] = 8'd71;
    sbox_0[23] = 8'd240;
    sbox_0[24] = 8'd173;
    sbox_0[25] = 8'd212;
    sbox_0[26] = 8'd162;
    sbox_0[27] = 8'd175;
    sbox_0[28] = 8'd156;
    sbox_0[29] = 8'd164;
    sbox_0[30] = 8'd114;
    sbox_0[31] = 8'd192;
    sbox_0[32] = 8'd183;
    sbox_0[33] = 8'd253;
    sbox_0[34] = 8'd147;
    sbox_0[35] = 8'd38;
    sbox_0[36] = 8'd54;
    sbox_0[37] = 8'd63;
    sbox_0[38] = 8'd247;
    sbox_0[39] = 8'd204;
    sbox_0[40] = 8'd52;
    sbox_0[41] = 8'd165;
    sbox_0[42] = 8'd229;
    sbox_0[43] = 8'd241;
    sbox_0[44] = 8'd113;
    sbox_0[45] = 8'd216;
    sbox_0[46] = 8'd49;
    sbox_0[47] = 8'd21;
    sbox_0[48] = 8'd4;
    sbox_0[49] = 8'd199;
    sbox_0[50] = 8'd35;
    sbox_0[51] = 8'd195;
    sbox_0[52] = 8'd24;
    sbox_0[53] = 8'd150;
    sbox_0[54] = 8'd5;
    sbox_0[55] = 8'd154;
    sbox_0[56] = 8'd7;
    sbox_0[57] = 8'd18;
    sbox_0[58] = 8'd128;
    sbox_0[59] = 8'd226;
    sbox_0[60] = 8'd235;
    sbox_0[61] = 8'd39;
    sbox_0[62] = 8'd178;
    sbox_0[63] = 8'd117;
    sbox_0[64] = 8'd9;
    sbox_0[65] = 8'd131;
    sbox_0[66] = 8'd44;
    sbox_0[67] = 8'd26;
    sbox_0[68] = 8'd27;
    sbox_0[69] = 8'd110;
    sbox_0[70] = 8'd90;
    sbox_0[71] = 8'd160;
    sbox_0[72] = 8'd82;
    sbox_0[73] = 8'd59;
    sbox_0[74] = 8'd214;
    sbox_0[75] = 8'd179;
    sbox_0[76] = 8'd41;
    sbox_0[77] = 8'd227;
    sbox_0[78] = 8'd47;
    sbox_0[79] = 8'd132;
    sbox_0[80] = 8'd83;
    sbox_0[81] = 8'd209;
    sbox_0[82] = 8'd0;
    sbox_0[83] = 8'd237;
    sbox_0[84] = 8'd32;
    sbox_0[85] = 8'd252;
    sbox_0[86] = 8'd177;
    sbox_0[87] = 8'd91;
    sbox_0[88] = 8'd106;
    sbox_0[89] = 8'd203;
    sbox_0[90] = 8'd190;
    sbox_0[91] = 8'd57;
    sbox_0[92] = 8'd74;
    sbox_0[93] = 8'd76;
    sbox_0[94] = 8'd88;
    sbox_0[95] = 8'd207;
    sbox_0[96] = 8'd208;
    sbox_0[97] = 8'd239;
    sbox_0[98] = 8'd170;
    sbox_0[99] = 8'd251;
    sbox_0[100] = 8'd67;
    sbox_0[101] = 8'd77;
    sbox_0[102] = 8'd51;
    sbox_0[103] = 8'd133;
    sbox_0[104] = 8'd69;
    sbox_0[105] = 8'd249;
    sbox_0[106] = 8'd2;
    sbox_0[107] = 8'd127;
    sbox_0[108] = 8'd80;
    sbox_0[109] = 8'd60;
    sbox_0[110] = 8'd159;
    sbox_0[111] = 8'd168;
    sbox_0[112] = 8'd81;
    sbox_0[113] = 8'd163;
    sbox_0[114] = 8'd64;
    sbox_0[115] = 8'd143;
    sbox_0[116] = 8'd146;
    sbox_0[117] = 8'd157;
    sbox_0[118] = 8'd56;
    sbox_0[119] = 8'd245;
    sbox_0[120] = 8'd188;
    sbox_0[121] = 8'd182;
    sbox_0[122] = 8'd218;
    sbox_0[123] = 8'd33;
    sbox_0[124] = 8'd16;
    sbox_0[125] = 8'd255;
    sbox_0[126] = 8'd243;
    sbox_0[127] = 8'd210;
    sbox_0[128] = 8'd205;
    sbox_0[129] = 8'd12;
    sbox_0[130] = 8'd19;
    sbox_0[131] = 8'd236;
    sbox_0[132] = 8'd95;
    sbox_0[133] = 8'd151;
    sbox_0[134] = 8'd68;
    sbox_0[135] = 8'd23;
    sbox_0[136] = 8'd196;
    sbox_0[137] = 8'd167;
    sbox_0[138] = 8'd126;
    sbox_0[139] = 8'd61;
    sbox_0[140] = 8'd100;
    sbox_0[141] = 8'd93;
    sbox_0[142] = 8'd25;
    sbox_0[143] = 8'd115;
    sbox_0[144] = 8'd96;
    sbox_0[145] = 8'd129;
    sbox_0[146] = 8'd79;
    sbox_0[147] = 8'd220;
    sbox_0[148] = 8'd34;
    sbox_0[149] = 8'd42;
    sbox_0[150] = 8'd144;
    sbox_0[151] = 8'd136;
    sbox_0[152] = 8'd70;
    sbox_0[153] = 8'd238;
    sbox_0[154] = 8'd184;
    sbox_0[155] = 8'd20;
    sbox_0[156] = 8'd222;
    sbox_0[157] = 8'd94;
    sbox_0[158] = 8'd11;
    sbox_0[159] = 8'd219;
    sbox_0[160] = 8'd224;
    sbox_0[161] = 8'd50;
    sbox_0[162] = 8'd58;
    sbox_0[163] = 8'd10;
    sbox_0[164] = 8'd73;
    sbox_0[165] = 8'd6;
    sbox_0[166] = 8'd36;
    sbox_0[167] = 8'd92;
    sbox_0[168] = 8'd194;
    sbox_0[169] = 8'd211;
    sbox_0[170] = 8'd172;
    sbox_0[171] = 8'd98;
    sbox_0[172] = 8'd145;
    sbox_0[173] = 8'd149;
    sbox_0[174] = 8'd228;
    sbox_0[175] = 8'd121;
    sbox_0[176] = 8'd231;
    sbox_0[177] = 8'd200;
    sbox_0[178] = 8'd55;
    sbox_0[179] = 8'd109;
    sbox_0[180] = 8'd141;
    sbox_0[181] = 8'd213;
    sbox_0[182] = 8'd78;
    sbox_0[183] = 8'd169;
    sbox_0[184] = 8'd108;
    sbox_0[185] = 8'd86;
    sbox_0[186] = 8'd244;
    sbox_0[187] = 8'd234;
    sbox_0[188] = 8'd101;
    sbox_0[189] = 8'd122;
    sbox_0[190] = 8'd174;
    sbox_0[191] = 8'd8;
    sbox_0[192] = 8'd186;
    sbox_0[193] = 8'd120;
    sbox_0[194] = 8'd37;
    sbox_0[195] = 8'd46;
    sbox_0[196] = 8'd28;
    sbox_0[197] = 8'd166;
    sbox_0[198] = 8'd180;
    sbox_0[199] = 8'd198;
    sbox_0[200] = 8'd232;
    sbox_0[201] = 8'd221;
    sbox_0[202] = 8'd116;
    sbox_0[203] = 8'd31;
    sbox_0[204] = 8'd75;
    sbox_0[205] = 8'd189;
    sbox_0[206] = 8'd139;
    sbox_0[207] = 8'd138;
    sbox_0[208] = 8'd112;
    sbox_0[209] = 8'd62;
    sbox_0[210] = 8'd181;
    sbox_0[211] = 8'd102;
    sbox_0[212] = 8'd72;
    sbox_0[213] = 8'd3;
    sbox_0[214] = 8'd246;
    sbox_0[215] = 8'd14;
    sbox_0[216] = 8'd97;
    sbox_0[217] = 8'd53;
    sbox_0[218] = 8'd87;
    sbox_0[219] = 8'd185;
    sbox_0[220] = 8'd134;
    sbox_0[221] = 8'd193;
    sbox_0[222] = 8'd29;
    sbox_0[223] = 8'd158;
    sbox_0[224] = 8'd225;
    sbox_0[225] = 8'd248;
    sbox_0[226] = 8'd152;
    sbox_0[227] = 8'd17;
    sbox_0[228] = 8'd105;
    sbox_0[229] = 8'd217;
    sbox_0[230] = 8'd142;
    sbox_0[231] = 8'd148;
    sbox_0[232] = 8'd155;
    sbox_0[233] = 8'd30;
    sbox_0[234] = 8'd135;
    sbox_0[235] = 8'd233;
    sbox_0[236] = 8'd206;
    sbox_0[237] = 8'd85;
    sbox_0[238] = 8'd40;
    sbox_0[239] = 8'd223;
    sbox_0[240] = 8'd140;
    sbox_0[241] = 8'd161;
    sbox_0[242] = 8'd137;
    sbox_0[243] = 8'd13;
    sbox_0[244] = 8'd191;
    sbox_0[245] = 8'd230;
    sbox_0[246] = 8'd66;
    sbox_0[247] = 8'd104;
    sbox_0[248] = 8'd65;
    sbox_0[249] = 8'd153;
    sbox_0[250] = 8'd45;
    sbox_0[251] = 8'd15;
    sbox_0[252] = 8'd176;
    sbox_0[253] = 8'd84;
    sbox_0[254] = 8'd187;
    sbox_0[255] = 8'd22;
    sbox_1[0] = 8'd99;
    sbox_1[1] = 8'd124;
    sbox_1[2] = 8'd119;
    sbox_1[3] = 8'd123;
    sbox_1[4] = 8'd242;
    sbox_1[5] = 8'd107;
    sbox_1[6] = 8'd111;
    sbox_1[7] = 8'd197;
    sbox_1[8] = 8'd48;
    sbox_1[9] = 8'd1;
    sbox_1[10] = 8'd103;
    sbox_1[11] = 8'd43;
    sbox_1[12] = 8'd254;
    sbox_1[13] = 8'd215;
    sbox_1[14] = 8'd171;
    sbox_1[15] = 8'd118;
    sbox_1[16] = 8'd202;
    sbox_1[17] = 8'd130;
    sbox_1[18] = 8'd201;
    sbox_1[19] = 8'd125;
    sbox_1[20] = 8'd250;
    sbox_1[21] = 8'd89;
    sbox_1[22] = 8'd71;
    sbox_1[23] = 8'd240;
    sbox_1[24] = 8'd173;
    sbox_1[25] = 8'd212;
    sbox_1[26] = 8'd162;
    sbox_1[27] = 8'd175;
    sbox_1[28] = 8'd156;
    sbox_1[29] = 8'd164;
    sbox_1[30] = 8'd114;
    sbox_1[31] = 8'd192;
    sbox_1[32] = 8'd183;
    sbox_1[33] = 8'd253;
    sbox_1[34] = 8'd147;
    sbox_1[35] = 8'd38;
    sbox_1[36] = 8'd54;
    sbox_1[37] = 8'd63;
    sbox_1[38] = 8'd247;
    sbox_1[39] = 8'd204;
    sbox_1[40] = 8'd52;
    sbox_1[41] = 8'd165;
    sbox_1[42] = 8'd229;
    sbox_1[43] = 8'd241;
    sbox_1[44] = 8'd113;
    sbox_1[45] = 8'd216;
    sbox_1[46] = 8'd49;
    sbox_1[47] = 8'd21;
    sbox_1[48] = 8'd4;
    sbox_1[49] = 8'd199;
    sbox_1[50] = 8'd35;
    sbox_1[51] = 8'd195;
    sbox_1[52] = 8'd24;
    sbox_1[53] = 8'd150;
    sbox_1[54] = 8'd5;
    sbox_1[55] = 8'd154;
    sbox_1[56] = 8'd7;
    sbox_1[57] = 8'd18;
    sbox_1[58] = 8'd128;
    sbox_1[59] = 8'd226;
    sbox_1[60] = 8'd235;
    sbox_1[61] = 8'd39;
    sbox_1[62] = 8'd178;
    sbox_1[63] = 8'd117;
    sbox_1[64] = 8'd9;
    sbox_1[65] = 8'd131;
    sbox_1[66] = 8'd44;
    sbox_1[67] = 8'd26;
    sbox_1[68] = 8'd27;
    sbox_1[69] = 8'd110;
    sbox_1[70] = 8'd90;
    sbox_1[71] = 8'd160;
    sbox_1[72] = 8'd82;
    sbox_1[73] = 8'd59;
    sbox_1[74] = 8'd214;
    sbox_1[75] = 8'd179;
    sbox_1[76] = 8'd41;
    sbox_1[77] = 8'd227;
    sbox_1[78] = 8'd47;
    sbox_1[79] = 8'd132;
    sbox_1[80] = 8'd83;
    sbox_1[81] = 8'd209;
    sbox_1[82] = 8'd0;
    sbox_1[83] = 8'd237;
    sbox_1[84] = 8'd32;
    sbox_1[85] = 8'd252;
    sbox_1[86] = 8'd177;
    sbox_1[87] = 8'd91;
    sbox_1[88] = 8'd106;
    sbox_1[89] = 8'd203;
    sbox_1[90] = 8'd190;
    sbox_1[91] = 8'd57;
    sbox_1[92] = 8'd74;
    sbox_1[93] = 8'd76;
    sbox_1[94] = 8'd88;
    sbox_1[95] = 8'd207;
    sbox_1[96] = 8'd208;
    sbox_1[97] = 8'd239;
    sbox_1[98] = 8'd170;
    sbox_1[99] = 8'd251;
    sbox_1[100] = 8'd67;
    sbox_1[101] = 8'd77;
    sbox_1[102] = 8'd51;
    sbox_1[103] = 8'd133;
    sbox_1[104] = 8'd69;
    sbox_1[105] = 8'd249;
    sbox_1[106] = 8'd2;
    sbox_1[107] = 8'd127;
    sbox_1[108] = 8'd80;
    sbox_1[109] = 8'd60;
    sbox_1[110] = 8'd159;
    sbox_1[111] = 8'd168;
    sbox_1[112] = 8'd81;
    sbox_1[113] = 8'd163;
    sbox_1[114] = 8'd64;
    sbox_1[115] = 8'd143;
    sbox_1[116] = 8'd146;
    sbox_1[117] = 8'd157;
    sbox_1[118] = 8'd56;
    sbox_1[119] = 8'd245;
    sbox_1[120] = 8'd188;
    sbox_1[121] = 8'd182;
    sbox_1[122] = 8'd218;
    sbox_1[123] = 8'd33;
    sbox_1[124] = 8'd16;
    sbox_1[125] = 8'd255;
    sbox_1[126] = 8'd243;
    sbox_1[127] = 8'd210;
    sbox_1[128] = 8'd205;
    sbox_1[129] = 8'd12;
    sbox_1[130] = 8'd19;
    sbox_1[131] = 8'd236;
    sbox_1[132] = 8'd95;
    sbox_1[133] = 8'd151;
    sbox_1[134] = 8'd68;
    sbox_1[135] = 8'd23;
    sbox_1[136] = 8'd196;
    sbox_1[137] = 8'd167;
    sbox_1[138] = 8'd126;
    sbox_1[139] = 8'd61;
    sbox_1[140] = 8'd100;
    sbox_1[141] = 8'd93;
    sbox_1[142] = 8'd25;
    sbox_1[143] = 8'd115;
    sbox_1[144] = 8'd96;
    sbox_1[145] = 8'd129;
    sbox_1[146] = 8'd79;
    sbox_1[147] = 8'd220;
    sbox_1[148] = 8'd34;
    sbox_1[149] = 8'd42;
    sbox_1[150] = 8'd144;
    sbox_1[151] = 8'd136;
    sbox_1[152] = 8'd70;
    sbox_1[153] = 8'd238;
    sbox_1[154] = 8'd184;
    sbox_1[155] = 8'd20;
    sbox_1[156] = 8'd222;
    sbox_1[157] = 8'd94;
    sbox_1[158] = 8'd11;
    sbox_1[159] = 8'd219;
    sbox_1[160] = 8'd224;
    sbox_1[161] = 8'd50;
    sbox_1[162] = 8'd58;
    sbox_1[163] = 8'd10;
    sbox_1[164] = 8'd73;
    sbox_1[165] = 8'd6;
    sbox_1[166] = 8'd36;
    sbox_1[167] = 8'd92;
    sbox_1[168] = 8'd194;
    sbox_1[169] = 8'd211;
    sbox_1[170] = 8'd172;
    sbox_1[171] = 8'd98;
    sbox_1[172] = 8'd145;
    sbox_1[173] = 8'd149;
    sbox_1[174] = 8'd228;
    sbox_1[175] = 8'd121;
    sbox_1[176] = 8'd231;
    sbox_1[177] = 8'd200;
    sbox_1[178] = 8'd55;
    sbox_1[179] = 8'd109;
    sbox_1[180] = 8'd141;
    sbox_1[181] = 8'd213;
    sbox_1[182] = 8'd78;
    sbox_1[183] = 8'd169;
    sbox_1[184] = 8'd108;
    sbox_1[185] = 8'd86;
    sbox_1[186] = 8'd244;
    sbox_1[187] = 8'd234;
    sbox_1[188] = 8'd101;
    sbox_1[189] = 8'd122;
    sbox_1[190] = 8'd174;
    sbox_1[191] = 8'd8;
    sbox_1[192] = 8'd186;
    sbox_1[193] = 8'd120;
    sbox_1[194] = 8'd37;
    sbox_1[195] = 8'd46;
    sbox_1[196] = 8'd28;
    sbox_1[197] = 8'd166;
    sbox_1[198] = 8'd180;
    sbox_1[199] = 8'd198;
    sbox_1[200] = 8'd232;
    sbox_1[201] = 8'd221;
    sbox_1[202] = 8'd116;
    sbox_1[203] = 8'd31;
    sbox_1[204] = 8'd75;
    sbox_1[205] = 8'd189;
    sbox_1[206] = 8'd139;
    sbox_1[207] = 8'd138;
    sbox_1[208] = 8'd112;
    sbox_1[209] = 8'd62;
    sbox_1[210] = 8'd181;
    sbox_1[211] = 8'd102;
    sbox_1[212] = 8'd72;
    sbox_1[213] = 8'd3;
    sbox_1[214] = 8'd246;
    sbox_1[215] = 8'd14;
    sbox_1[216] = 8'd97;
    sbox_1[217] = 8'd53;
    sbox_1[218] = 8'd87;
    sbox_1[219] = 8'd185;
    sbox_1[220] = 8'd134;
    sbox_1[221] = 8'd193;
    sbox_1[222] = 8'd29;
    sbox_1[223] = 8'd158;
    sbox_1[224] = 8'd225;
    sbox_1[225] = 8'd248;
    sbox_1[226] = 8'd152;
    sbox_1[227] = 8'd17;
    sbox_1[228] = 8'd105;
    sbox_1[229] = 8'd217;
    sbox_1[230] = 8'd142;
    sbox_1[231] = 8'd148;
    sbox_1[232] = 8'd155;
    sbox_1[233] = 8'd30;
    sbox_1[234] = 8'd135;
    sbox_1[235] = 8'd233;
    sbox_1[236] = 8'd206;
    sbox_1[237] = 8'd85;
    sbox_1[238] = 8'd40;
    sbox_1[239] = 8'd223;
    sbox_1[240] = 8'd140;
    sbox_1[241] = 8'd161;
    sbox_1[242] = 8'd137;
    sbox_1[243] = 8'd13;
    sbox_1[244] = 8'd191;
    sbox_1[245] = 8'd230;
    sbox_1[246] = 8'd66;
    sbox_1[247] = 8'd104;
    sbox_1[248] = 8'd65;
    sbox_1[249] = 8'd153;
    sbox_1[250] = 8'd45;
    sbox_1[251] = 8'd15;
    sbox_1[252] = 8'd176;
    sbox_1[253] = 8'd84;
    sbox_1[254] = 8'd187;
    sbox_1[255] = 8'd22;
    sbox_2[0] = 8'd99;
    sbox_2[1] = 8'd124;
    sbox_2[2] = 8'd119;
    sbox_2[3] = 8'd123;
    sbox_2[4] = 8'd242;
    sbox_2[5] = 8'd107;
    sbox_2[6] = 8'd111;
    sbox_2[7] = 8'd197;
    sbox_2[8] = 8'd48;
    sbox_2[9] = 8'd1;
    sbox_2[10] = 8'd103;
    sbox_2[11] = 8'd43;
    sbox_2[12] = 8'd254;
    sbox_2[13] = 8'd215;
    sbox_2[14] = 8'd171;
    sbox_2[15] = 8'd118;
    sbox_2[16] = 8'd202;
    sbox_2[17] = 8'd130;
    sbox_2[18] = 8'd201;
    sbox_2[19] = 8'd125;
    sbox_2[20] = 8'd250;
    sbox_2[21] = 8'd89;
    sbox_2[22] = 8'd71;
    sbox_2[23] = 8'd240;
    sbox_2[24] = 8'd173;
    sbox_2[25] = 8'd212;
    sbox_2[26] = 8'd162;
    sbox_2[27] = 8'd175;
    sbox_2[28] = 8'd156;
    sbox_2[29] = 8'd164;
    sbox_2[30] = 8'd114;
    sbox_2[31] = 8'd192;
    sbox_2[32] = 8'd183;
    sbox_2[33] = 8'd253;
    sbox_2[34] = 8'd147;
    sbox_2[35] = 8'd38;
    sbox_2[36] = 8'd54;
    sbox_2[37] = 8'd63;
    sbox_2[38] = 8'd247;
    sbox_2[39] = 8'd204;
    sbox_2[40] = 8'd52;
    sbox_2[41] = 8'd165;
    sbox_2[42] = 8'd229;
    sbox_2[43] = 8'd241;
    sbox_2[44] = 8'd113;
    sbox_2[45] = 8'd216;
    sbox_2[46] = 8'd49;
    sbox_2[47] = 8'd21;
    sbox_2[48] = 8'd4;
    sbox_2[49] = 8'd199;
    sbox_2[50] = 8'd35;
    sbox_2[51] = 8'd195;
    sbox_2[52] = 8'd24;
    sbox_2[53] = 8'd150;
    sbox_2[54] = 8'd5;
    sbox_2[55] = 8'd154;
    sbox_2[56] = 8'd7;
    sbox_2[57] = 8'd18;
    sbox_2[58] = 8'd128;
    sbox_2[59] = 8'd226;
    sbox_2[60] = 8'd235;
    sbox_2[61] = 8'd39;
    sbox_2[62] = 8'd178;
    sbox_2[63] = 8'd117;
    sbox_2[64] = 8'd9;
    sbox_2[65] = 8'd131;
    sbox_2[66] = 8'd44;
    sbox_2[67] = 8'd26;
    sbox_2[68] = 8'd27;
    sbox_2[69] = 8'd110;
    sbox_2[70] = 8'd90;
    sbox_2[71] = 8'd160;
    sbox_2[72] = 8'd82;
    sbox_2[73] = 8'd59;
    sbox_2[74] = 8'd214;
    sbox_2[75] = 8'd179;
    sbox_2[76] = 8'd41;
    sbox_2[77] = 8'd227;
    sbox_2[78] = 8'd47;
    sbox_2[79] = 8'd132;
    sbox_2[80] = 8'd83;
    sbox_2[81] = 8'd209;
    sbox_2[82] = 8'd0;
    sbox_2[83] = 8'd237;
    sbox_2[84] = 8'd32;
    sbox_2[85] = 8'd252;
    sbox_2[86] = 8'd177;
    sbox_2[87] = 8'd91;
    sbox_2[88] = 8'd106;
    sbox_2[89] = 8'd203;
    sbox_2[90] = 8'd190;
    sbox_2[91] = 8'd57;
    sbox_2[92] = 8'd74;
    sbox_2[93] = 8'd76;
    sbox_2[94] = 8'd88;
    sbox_2[95] = 8'd207;
    sbox_2[96] = 8'd208;
    sbox_2[97] = 8'd239;
    sbox_2[98] = 8'd170;
    sbox_2[99] = 8'd251;
    sbox_2[100] = 8'd67;
    sbox_2[101] = 8'd77;
    sbox_2[102] = 8'd51;
    sbox_2[103] = 8'd133;
    sbox_2[104] = 8'd69;
    sbox_2[105] = 8'd249;
    sbox_2[106] = 8'd2;
    sbox_2[107] = 8'd127;
    sbox_2[108] = 8'd80;
    sbox_2[109] = 8'd60;
    sbox_2[110] = 8'd159;
    sbox_2[111] = 8'd168;
    sbox_2[112] = 8'd81;
    sbox_2[113] = 8'd163;
    sbox_2[114] = 8'd64;
    sbox_2[115] = 8'd143;
    sbox_2[116] = 8'd146;
    sbox_2[117] = 8'd157;
    sbox_2[118] = 8'd56;
    sbox_2[119] = 8'd245;
    sbox_2[120] = 8'd188;
    sbox_2[121] = 8'd182;
    sbox_2[122] = 8'd218;
    sbox_2[123] = 8'd33;
    sbox_2[124] = 8'd16;
    sbox_2[125] = 8'd255;
    sbox_2[126] = 8'd243;
    sbox_2[127] = 8'd210;
    sbox_2[128] = 8'd205;
    sbox_2[129] = 8'd12;
    sbox_2[130] = 8'd19;
    sbox_2[131] = 8'd236;
    sbox_2[132] = 8'd95;
    sbox_2[133] = 8'd151;
    sbox_2[134] = 8'd68;
    sbox_2[135] = 8'd23;
    sbox_2[136] = 8'd196;
    sbox_2[137] = 8'd167;
    sbox_2[138] = 8'd126;
    sbox_2[139] = 8'd61;
    sbox_2[140] = 8'd100;
    sbox_2[141] = 8'd93;
    sbox_2[142] = 8'd25;
    sbox_2[143] = 8'd115;
    sbox_2[144] = 8'd96;
    sbox_2[145] = 8'd129;
    sbox_2[146] = 8'd79;
    sbox_2[147] = 8'd220;
    sbox_2[148] = 8'd34;
    sbox_2[149] = 8'd42;
    sbox_2[150] = 8'd144;
    sbox_2[151] = 8'd136;
    sbox_2[152] = 8'd70;
    sbox_2[153] = 8'd238;
    sbox_2[154] = 8'd184;
    sbox_2[155] = 8'd20;
    sbox_2[156] = 8'd222;
    sbox_2[157] = 8'd94;
    sbox_2[158] = 8'd11;
    sbox_2[159] = 8'd219;
    sbox_2[160] = 8'd224;
    sbox_2[161] = 8'd50;
    sbox_2[162] = 8'd58;
    sbox_2[163] = 8'd10;
    sbox_2[164] = 8'd73;
    sbox_2[165] = 8'd6;
    sbox_2[166] = 8'd36;
    sbox_2[167] = 8'd92;
    sbox_2[168] = 8'd194;
    sbox_2[169] = 8'd211;
    sbox_2[170] = 8'd172;
    sbox_2[171] = 8'd98;
    sbox_2[172] = 8'd145;
    sbox_2[173] = 8'd149;
    sbox_2[174] = 8'd228;
    sbox_2[175] = 8'd121;
    sbox_2[176] = 8'd231;
    sbox_2[177] = 8'd200;
    sbox_2[178] = 8'd55;
    sbox_2[179] = 8'd109;
    sbox_2[180] = 8'd141;
    sbox_2[181] = 8'd213;
    sbox_2[182] = 8'd78;
    sbox_2[183] = 8'd169;
    sbox_2[184] = 8'd108;
    sbox_2[185] = 8'd86;
    sbox_2[186] = 8'd244;
    sbox_2[187] = 8'd234;
    sbox_2[188] = 8'd101;
    sbox_2[189] = 8'd122;
    sbox_2[190] = 8'd174;
    sbox_2[191] = 8'd8;
    sbox_2[192] = 8'd186;
    sbox_2[193] = 8'd120;
    sbox_2[194] = 8'd37;
    sbox_2[195] = 8'd46;
    sbox_2[196] = 8'd28;
    sbox_2[197] = 8'd166;
    sbox_2[198] = 8'd180;
    sbox_2[199] = 8'd198;
    sbox_2[200] = 8'd232;
    sbox_2[201] = 8'd221;
    sbox_2[202] = 8'd116;
    sbox_2[203] = 8'd31;
    sbox_2[204] = 8'd75;
    sbox_2[205] = 8'd189;
    sbox_2[206] = 8'd139;
    sbox_2[207] = 8'd138;
    sbox_2[208] = 8'd112;
    sbox_2[209] = 8'd62;
    sbox_2[210] = 8'd181;
    sbox_2[211] = 8'd102;
    sbox_2[212] = 8'd72;
    sbox_2[213] = 8'd3;
    sbox_2[214] = 8'd246;
    sbox_2[215] = 8'd14;
    sbox_2[216] = 8'd97;
    sbox_2[217] = 8'd53;
    sbox_2[218] = 8'd87;
    sbox_2[219] = 8'd185;
    sbox_2[220] = 8'd134;
    sbox_2[221] = 8'd193;
    sbox_2[222] = 8'd29;
    sbox_2[223] = 8'd158;
    sbox_2[224] = 8'd225;
    sbox_2[225] = 8'd248;
    sbox_2[226] = 8'd152;
    sbox_2[227] = 8'd17;
    sbox_2[228] = 8'd105;
    sbox_2[229] = 8'd217;
    sbox_2[230] = 8'd142;
    sbox_2[231] = 8'd148;
    sbox_2[232] = 8'd155;
    sbox_2[233] = 8'd30;
    sbox_2[234] = 8'd135;
    sbox_2[235] = 8'd233;
    sbox_2[236] = 8'd206;
    sbox_2[237] = 8'd85;
    sbox_2[238] = 8'd40;
    sbox_2[239] = 8'd223;
    sbox_2[240] = 8'd140;
    sbox_2[241] = 8'd161;
    sbox_2[242] = 8'd137;
    sbox_2[243] = 8'd13;
    sbox_2[244] = 8'd191;
    sbox_2[245] = 8'd230;
    sbox_2[246] = 8'd66;
    sbox_2[247] = 8'd104;
    sbox_2[248] = 8'd65;
    sbox_2[249] = 8'd153;
    sbox_2[250] = 8'd45;
    sbox_2[251] = 8'd15;
    sbox_2[252] = 8'd176;
    sbox_2[253] = 8'd84;
    sbox_2[254] = 8'd187;
    sbox_2[255] = 8'd22;
    sbox_3[0] = 8'd99;
    sbox_3[1] = 8'd124;
    sbox_3[2] = 8'd119;
    sbox_3[3] = 8'd123;
    sbox_3[4] = 8'd242;
    sbox_3[5] = 8'd107;
    sbox_3[6] = 8'd111;
    sbox_3[7] = 8'd197;
    sbox_3[8] = 8'd48;
    sbox_3[9] = 8'd1;
    sbox_3[10] = 8'd103;
    sbox_3[11] = 8'd43;
    sbox_3[12] = 8'd254;
    sbox_3[13] = 8'd215;
    sbox_3[14] = 8'd171;
    sbox_3[15] = 8'd118;
    sbox_3[16] = 8'd202;
    sbox_3[17] = 8'd130;
    sbox_3[18] = 8'd201;
    sbox_3[19] = 8'd125;
    sbox_3[20] = 8'd250;
    sbox_3[21] = 8'd89;
    sbox_3[22] = 8'd71;
    sbox_3[23] = 8'd240;
    sbox_3[24] = 8'd173;
    sbox_3[25] = 8'd212;
    sbox_3[26] = 8'd162;
    sbox_3[27] = 8'd175;
    sbox_3[28] = 8'd156;
    sbox_3[29] = 8'd164;
    sbox_3[30] = 8'd114;
    sbox_3[31] = 8'd192;
    sbox_3[32] = 8'd183;
    sbox_3[33] = 8'd253;
    sbox_3[34] = 8'd147;
    sbox_3[35] = 8'd38;
    sbox_3[36] = 8'd54;
    sbox_3[37] = 8'd63;
    sbox_3[38] = 8'd247;
    sbox_3[39] = 8'd204;
    sbox_3[40] = 8'd52;
    sbox_3[41] = 8'd165;
    sbox_3[42] = 8'd229;
    sbox_3[43] = 8'd241;
    sbox_3[44] = 8'd113;
    sbox_3[45] = 8'd216;
    sbox_3[46] = 8'd49;
    sbox_3[47] = 8'd21;
    sbox_3[48] = 8'd4;
    sbox_3[49] = 8'd199;
    sbox_3[50] = 8'd35;
    sbox_3[51] = 8'd195;
    sbox_3[52] = 8'd24;
    sbox_3[53] = 8'd150;
    sbox_3[54] = 8'd5;
    sbox_3[55] = 8'd154;
    sbox_3[56] = 8'd7;
    sbox_3[57] = 8'd18;
    sbox_3[58] = 8'd128;
    sbox_3[59] = 8'd226;
    sbox_3[60] = 8'd235;
    sbox_3[61] = 8'd39;
    sbox_3[62] = 8'd178;
    sbox_3[63] = 8'd117;
    sbox_3[64] = 8'd9;
    sbox_3[65] = 8'd131;
    sbox_3[66] = 8'd44;
    sbox_3[67] = 8'd26;
    sbox_3[68] = 8'd27;
    sbox_3[69] = 8'd110;
    sbox_3[70] = 8'd90;
    sbox_3[71] = 8'd160;
    sbox_3[72] = 8'd82;
    sbox_3[73] = 8'd59;
    sbox_3[74] = 8'd214;
    sbox_3[75] = 8'd179;
    sbox_3[76] = 8'd41;
    sbox_3[77] = 8'd227;
    sbox_3[78] = 8'd47;
    sbox_3[79] = 8'd132;
    sbox_3[80] = 8'd83;
    sbox_3[81] = 8'd209;
    sbox_3[82] = 8'd0;
    sbox_3[83] = 8'd237;
    sbox_3[84] = 8'd32;
    sbox_3[85] = 8'd252;
    sbox_3[86] = 8'd177;
    sbox_3[87] = 8'd91;
    sbox_3[88] = 8'd106;
    sbox_3[89] = 8'd203;
    sbox_3[90] = 8'd190;
    sbox_3[91] = 8'd57;
    sbox_3[92] = 8'd74;
    sbox_3[93] = 8'd76;
    sbox_3[94] = 8'd88;
    sbox_3[95] = 8'd207;
    sbox_3[96] = 8'd208;
    sbox_3[97] = 8'd239;
    sbox_3[98] = 8'd170;
    sbox_3[99] = 8'd251;
    sbox_3[100] = 8'd67;
    sbox_3[101] = 8'd77;
    sbox_3[102] = 8'd51;
    sbox_3[103] = 8'd133;
    sbox_3[104] = 8'd69;
    sbox_3[105] = 8'd249;
    sbox_3[106] = 8'd2;
    sbox_3[107] = 8'd127;
    sbox_3[108] = 8'd80;
    sbox_3[109] = 8'd60;
    sbox_3[110] = 8'd159;
    sbox_3[111] = 8'd168;
    sbox_3[112] = 8'd81;
    sbox_3[113] = 8'd163;
    sbox_3[114] = 8'd64;
    sbox_3[115] = 8'd143;
    sbox_3[116] = 8'd146;
    sbox_3[117] = 8'd157;
    sbox_3[118] = 8'd56;
    sbox_3[119] = 8'd245;
    sbox_3[120] = 8'd188;
    sbox_3[121] = 8'd182;
    sbox_3[122] = 8'd218;
    sbox_3[123] = 8'd33;
    sbox_3[124] = 8'd16;
    sbox_3[125] = 8'd255;
    sbox_3[126] = 8'd243;
    sbox_3[127] = 8'd210;
    sbox_3[128] = 8'd205;
    sbox_3[129] = 8'd12;
    sbox_3[130] = 8'd19;
    sbox_3[131] = 8'd236;
    sbox_3[132] = 8'd95;
    sbox_3[133] = 8'd151;
    sbox_3[134] = 8'd68;
    sbox_3[135] = 8'd23;
    sbox_3[136] = 8'd196;
    sbox_3[137] = 8'd167;
    sbox_3[138] = 8'd126;
    sbox_3[139] = 8'd61;
    sbox_3[140] = 8'd100;
    sbox_3[141] = 8'd93;
    sbox_3[142] = 8'd25;
    sbox_3[143] = 8'd115;
    sbox_3[144] = 8'd96;
    sbox_3[145] = 8'd129;
    sbox_3[146] = 8'd79;
    sbox_3[147] = 8'd220;
    sbox_3[148] = 8'd34;
    sbox_3[149] = 8'd42;
    sbox_3[150] = 8'd144;
    sbox_3[151] = 8'd136;
    sbox_3[152] = 8'd70;
    sbox_3[153] = 8'd238;
    sbox_3[154] = 8'd184;
    sbox_3[155] = 8'd20;
    sbox_3[156] = 8'd222;
    sbox_3[157] = 8'd94;
    sbox_3[158] = 8'd11;
    sbox_3[159] = 8'd219;
    sbox_3[160] = 8'd224;
    sbox_3[161] = 8'd50;
    sbox_3[162] = 8'd58;
    sbox_3[163] = 8'd10;
    sbox_3[164] = 8'd73;
    sbox_3[165] = 8'd6;
    sbox_3[166] = 8'd36;
    sbox_3[167] = 8'd92;
    sbox_3[168] = 8'd194;
    sbox_3[169] = 8'd211;
    sbox_3[170] = 8'd172;
    sbox_3[171] = 8'd98;
    sbox_3[172] = 8'd145;
    sbox_3[173] = 8'd149;
    sbox_3[174] = 8'd228;
    sbox_3[175] = 8'd121;
    sbox_3[176] = 8'd231;
    sbox_3[177] = 8'd200;
    sbox_3[178] = 8'd55;
    sbox_3[179] = 8'd109;
    sbox_3[180] = 8'd141;
    sbox_3[181] = 8'd213;
    sbox_3[182] = 8'd78;
    sbox_3[183] = 8'd169;
    sbox_3[184] = 8'd108;
    sbox_3[185] = 8'd86;
    sbox_3[186] = 8'd244;
    sbox_3[187] = 8'd234;
    sbox_3[188] = 8'd101;
    sbox_3[189] = 8'd122;
    sbox_3[190] = 8'd174;
    sbox_3[191] = 8'd8;
    sbox_3[192] = 8'd186;
    sbox_3[193] = 8'd120;
    sbox_3[194] = 8'd37;
    sbox_3[195] = 8'd46;
    sbox_3[196] = 8'd28;
    sbox_3[197] = 8'd166;
    sbox_3[198] = 8'd180;
    sbox_3[199] = 8'd198;
    sbox_3[200] = 8'd232;
    sbox_3[201] = 8'd221;
    sbox_3[202] = 8'd116;
    sbox_3[203] = 8'd31;
    sbox_3[204] = 8'd75;
    sbox_3[205] = 8'd189;
    sbox_3[206] = 8'd139;
    sbox_3[207] = 8'd138;
    sbox_3[208] = 8'd112;
    sbox_3[209] = 8'd62;
    sbox_3[210] = 8'd181;
    sbox_3[211] = 8'd102;
    sbox_3[212] = 8'd72;
    sbox_3[213] = 8'd3;
    sbox_3[214] = 8'd246;
    sbox_3[215] = 8'd14;
    sbox_3[216] = 8'd97;
    sbox_3[217] = 8'd53;
    sbox_3[218] = 8'd87;
    sbox_3[219] = 8'd185;
    sbox_3[220] = 8'd134;
    sbox_3[221] = 8'd193;
    sbox_3[222] = 8'd29;
    sbox_3[223] = 8'd158;
    sbox_3[224] = 8'd225;
    sbox_3[225] = 8'd248;
    sbox_3[226] = 8'd152;
    sbox_3[227] = 8'd17;
    sbox_3[228] = 8'd105;
    sbox_3[229] = 8'd217;
    sbox_3[230] = 8'd142;
    sbox_3[231] = 8'd148;
    sbox_3[232] = 8'd155;
    sbox_3[233] = 8'd30;
    sbox_3[234] = 8'd135;
    sbox_3[235] = 8'd233;
    sbox_3[236] = 8'd206;
    sbox_3[237] = 8'd85;
    sbox_3[238] = 8'd40;
    sbox_3[239] = 8'd223;
    sbox_3[240] = 8'd140;
    sbox_3[241] = 8'd161;
    sbox_3[242] = 8'd137;
    sbox_3[243] = 8'd13;
    sbox_3[244] = 8'd191;
    sbox_3[245] = 8'd230;
    sbox_3[246] = 8'd66;
    sbox_3[247] = 8'd104;
    sbox_3[248] = 8'd65;
    sbox_3[249] = 8'd153;
    sbox_3[250] = 8'd45;
    sbox_3[251] = 8'd15;
    sbox_3[252] = 8'd176;
    sbox_3[253] = 8'd84;
    sbox_3[254] = 8'd187;
    sbox_3[255] = 8'd22;
    sbox_4[0] = 8'd99;
    sbox_4[1] = 8'd124;
    sbox_4[2] = 8'd119;
    sbox_4[3] = 8'd123;
    sbox_4[4] = 8'd242;
    sbox_4[5] = 8'd107;
    sbox_4[6] = 8'd111;
    sbox_4[7] = 8'd197;
    sbox_4[8] = 8'd48;
    sbox_4[9] = 8'd1;
    sbox_4[10] = 8'd103;
    sbox_4[11] = 8'd43;
    sbox_4[12] = 8'd254;
    sbox_4[13] = 8'd215;
    sbox_4[14] = 8'd171;
    sbox_4[15] = 8'd118;
    sbox_4[16] = 8'd202;
    sbox_4[17] = 8'd130;
    sbox_4[18] = 8'd201;
    sbox_4[19] = 8'd125;
    sbox_4[20] = 8'd250;
    sbox_4[21] = 8'd89;
    sbox_4[22] = 8'd71;
    sbox_4[23] = 8'd240;
    sbox_4[24] = 8'd173;
    sbox_4[25] = 8'd212;
    sbox_4[26] = 8'd162;
    sbox_4[27] = 8'd175;
    sbox_4[28] = 8'd156;
    sbox_4[29] = 8'd164;
    sbox_4[30] = 8'd114;
    sbox_4[31] = 8'd192;
    sbox_4[32] = 8'd183;
    sbox_4[33] = 8'd253;
    sbox_4[34] = 8'd147;
    sbox_4[35] = 8'd38;
    sbox_4[36] = 8'd54;
    sbox_4[37] = 8'd63;
    sbox_4[38] = 8'd247;
    sbox_4[39] = 8'd204;
    sbox_4[40] = 8'd52;
    sbox_4[41] = 8'd165;
    sbox_4[42] = 8'd229;
    sbox_4[43] = 8'd241;
    sbox_4[44] = 8'd113;
    sbox_4[45] = 8'd216;
    sbox_4[46] = 8'd49;
    sbox_4[47] = 8'd21;
    sbox_4[48] = 8'd4;
    sbox_4[49] = 8'd199;
    sbox_4[50] = 8'd35;
    sbox_4[51] = 8'd195;
    sbox_4[52] = 8'd24;
    sbox_4[53] = 8'd150;
    sbox_4[54] = 8'd5;
    sbox_4[55] = 8'd154;
    sbox_4[56] = 8'd7;
    sbox_4[57] = 8'd18;
    sbox_4[58] = 8'd128;
    sbox_4[59] = 8'd226;
    sbox_4[60] = 8'd235;
    sbox_4[61] = 8'd39;
    sbox_4[62] = 8'd178;
    sbox_4[63] = 8'd117;
    sbox_4[64] = 8'd9;
    sbox_4[65] = 8'd131;
    sbox_4[66] = 8'd44;
    sbox_4[67] = 8'd26;
    sbox_4[68] = 8'd27;
    sbox_4[69] = 8'd110;
    sbox_4[70] = 8'd90;
    sbox_4[71] = 8'd160;
    sbox_4[72] = 8'd82;
    sbox_4[73] = 8'd59;
    sbox_4[74] = 8'd214;
    sbox_4[75] = 8'd179;
    sbox_4[76] = 8'd41;
    sbox_4[77] = 8'd227;
    sbox_4[78] = 8'd47;
    sbox_4[79] = 8'd132;
    sbox_4[80] = 8'd83;
    sbox_4[81] = 8'd209;
    sbox_4[82] = 8'd0;
    sbox_4[83] = 8'd237;
    sbox_4[84] = 8'd32;
    sbox_4[85] = 8'd252;
    sbox_4[86] = 8'd177;
    sbox_4[87] = 8'd91;
    sbox_4[88] = 8'd106;
    sbox_4[89] = 8'd203;
    sbox_4[90] = 8'd190;
    sbox_4[91] = 8'd57;
    sbox_4[92] = 8'd74;
    sbox_4[93] = 8'd76;
    sbox_4[94] = 8'd88;
    sbox_4[95] = 8'd207;
    sbox_4[96] = 8'd208;
    sbox_4[97] = 8'd239;
    sbox_4[98] = 8'd170;
    sbox_4[99] = 8'd251;
    sbox_4[100] = 8'd67;
    sbox_4[101] = 8'd77;
    sbox_4[102] = 8'd51;
    sbox_4[103] = 8'd133;
    sbox_4[104] = 8'd69;
    sbox_4[105] = 8'd249;
    sbox_4[106] = 8'd2;
    sbox_4[107] = 8'd127;
    sbox_4[108] = 8'd80;
    sbox_4[109] = 8'd60;
    sbox_4[110] = 8'd159;
    sbox_4[111] = 8'd168;
    sbox_4[112] = 8'd81;
    sbox_4[113] = 8'd163;
    sbox_4[114] = 8'd64;
    sbox_4[115] = 8'd143;
    sbox_4[116] = 8'd146;
    sbox_4[117] = 8'd157;
    sbox_4[118] = 8'd56;
    sbox_4[119] = 8'd245;
    sbox_4[120] = 8'd188;
    sbox_4[121] = 8'd182;
    sbox_4[122] = 8'd218;
    sbox_4[123] = 8'd33;
    sbox_4[124] = 8'd16;
    sbox_4[125] = 8'd255;
    sbox_4[126] = 8'd243;
    sbox_4[127] = 8'd210;
    sbox_4[128] = 8'd205;
    sbox_4[129] = 8'd12;
    sbox_4[130] = 8'd19;
    sbox_4[131] = 8'd236;
    sbox_4[132] = 8'd95;
    sbox_4[133] = 8'd151;
    sbox_4[134] = 8'd68;
    sbox_4[135] = 8'd23;
    sbox_4[136] = 8'd196;
    sbox_4[137] = 8'd167;
    sbox_4[138] = 8'd126;
    sbox_4[139] = 8'd61;
    sbox_4[140] = 8'd100;
    sbox_4[141] = 8'd93;
    sbox_4[142] = 8'd25;
    sbox_4[143] = 8'd115;
    sbox_4[144] = 8'd96;
    sbox_4[145] = 8'd129;
    sbox_4[146] = 8'd79;
    sbox_4[147] = 8'd220;
    sbox_4[148] = 8'd34;
    sbox_4[149] = 8'd42;
    sbox_4[150] = 8'd144;
    sbox_4[151] = 8'd136;
    sbox_4[152] = 8'd70;
    sbox_4[153] = 8'd238;
    sbox_4[154] = 8'd184;
    sbox_4[155] = 8'd20;
    sbox_4[156] = 8'd222;
    sbox_4[157] = 8'd94;
    sbox_4[158] = 8'd11;
    sbox_4[159] = 8'd219;
    sbox_4[160] = 8'd224;
    sbox_4[161] = 8'd50;
    sbox_4[162] = 8'd58;
    sbox_4[163] = 8'd10;
    sbox_4[164] = 8'd73;
    sbox_4[165] = 8'd6;
    sbox_4[166] = 8'd36;
    sbox_4[167] = 8'd92;
    sbox_4[168] = 8'd194;
    sbox_4[169] = 8'd211;
    sbox_4[170] = 8'd172;
    sbox_4[171] = 8'd98;
    sbox_4[172] = 8'd145;
    sbox_4[173] = 8'd149;
    sbox_4[174] = 8'd228;
    sbox_4[175] = 8'd121;
    sbox_4[176] = 8'd231;
    sbox_4[177] = 8'd200;
    sbox_4[178] = 8'd55;
    sbox_4[179] = 8'd109;
    sbox_4[180] = 8'd141;
    sbox_4[181] = 8'd213;
    sbox_4[182] = 8'd78;
    sbox_4[183] = 8'd169;
    sbox_4[184] = 8'd108;
    sbox_4[185] = 8'd86;
    sbox_4[186] = 8'd244;
    sbox_4[187] = 8'd234;
    sbox_4[188] = 8'd101;
    sbox_4[189] = 8'd122;
    sbox_4[190] = 8'd174;
    sbox_4[191] = 8'd8;
    sbox_4[192] = 8'd186;
    sbox_4[193] = 8'd120;
    sbox_4[194] = 8'd37;
    sbox_4[195] = 8'd46;
    sbox_4[196] = 8'd28;
    sbox_4[197] = 8'd166;
    sbox_4[198] = 8'd180;
    sbox_4[199] = 8'd198;
    sbox_4[200] = 8'd232;
    sbox_4[201] = 8'd221;
    sbox_4[202] = 8'd116;
    sbox_4[203] = 8'd31;
    sbox_4[204] = 8'd75;
    sbox_4[205] = 8'd189;
    sbox_4[206] = 8'd139;
    sbox_4[207] = 8'd138;
    sbox_4[208] = 8'd112;
    sbox_4[209] = 8'd62;
    sbox_4[210] = 8'd181;
    sbox_4[211] = 8'd102;
    sbox_4[212] = 8'd72;
    sbox_4[213] = 8'd3;
    sbox_4[214] = 8'd246;
    sbox_4[215] = 8'd14;
    sbox_4[216] = 8'd97;
    sbox_4[217] = 8'd53;
    sbox_4[218] = 8'd87;
    sbox_4[219] = 8'd185;
    sbox_4[220] = 8'd134;
    sbox_4[221] = 8'd193;
    sbox_4[222] = 8'd29;
    sbox_4[223] = 8'd158;
    sbox_4[224] = 8'd225;
    sbox_4[225] = 8'd248;
    sbox_4[226] = 8'd152;
    sbox_4[227] = 8'd17;
    sbox_4[228] = 8'd105;
    sbox_4[229] = 8'd217;
    sbox_4[230] = 8'd142;
    sbox_4[231] = 8'd148;
    sbox_4[232] = 8'd155;
    sbox_4[233] = 8'd30;
    sbox_4[234] = 8'd135;
    sbox_4[235] = 8'd233;
    sbox_4[236] = 8'd206;
    sbox_4[237] = 8'd85;
    sbox_4[238] = 8'd40;
    sbox_4[239] = 8'd223;
    sbox_4[240] = 8'd140;
    sbox_4[241] = 8'd161;
    sbox_4[242] = 8'd137;
    sbox_4[243] = 8'd13;
    sbox_4[244] = 8'd191;
    sbox_4[245] = 8'd230;
    sbox_4[246] = 8'd66;
    sbox_4[247] = 8'd104;
    sbox_4[248] = 8'd65;
    sbox_4[249] = 8'd153;
    sbox_4[250] = 8'd45;
    sbox_4[251] = 8'd15;
    sbox_4[252] = 8'd176;
    sbox_4[253] = 8'd84;
    sbox_4[254] = 8'd187;
    sbox_4[255] = 8'd22;
    sbox_5[0] = 8'd99;
    sbox_5[1] = 8'd124;
    sbox_5[2] = 8'd119;
    sbox_5[3] = 8'd123;
    sbox_5[4] = 8'd242;
    sbox_5[5] = 8'd107;
    sbox_5[6] = 8'd111;
    sbox_5[7] = 8'd197;
    sbox_5[8] = 8'd48;
    sbox_5[9] = 8'd1;
    sbox_5[10] = 8'd103;
    sbox_5[11] = 8'd43;
    sbox_5[12] = 8'd254;
    sbox_5[13] = 8'd215;
    sbox_5[14] = 8'd171;
    sbox_5[15] = 8'd118;
    sbox_5[16] = 8'd202;
    sbox_5[17] = 8'd130;
    sbox_5[18] = 8'd201;
    sbox_5[19] = 8'd125;
    sbox_5[20] = 8'd250;
    sbox_5[21] = 8'd89;
    sbox_5[22] = 8'd71;
    sbox_5[23] = 8'd240;
    sbox_5[24] = 8'd173;
    sbox_5[25] = 8'd212;
    sbox_5[26] = 8'd162;
    sbox_5[27] = 8'd175;
    sbox_5[28] = 8'd156;
    sbox_5[29] = 8'd164;
    sbox_5[30] = 8'd114;
    sbox_5[31] = 8'd192;
    sbox_5[32] = 8'd183;
    sbox_5[33] = 8'd253;
    sbox_5[34] = 8'd147;
    sbox_5[35] = 8'd38;
    sbox_5[36] = 8'd54;
    sbox_5[37] = 8'd63;
    sbox_5[38] = 8'd247;
    sbox_5[39] = 8'd204;
    sbox_5[40] = 8'd52;
    sbox_5[41] = 8'd165;
    sbox_5[42] = 8'd229;
    sbox_5[43] = 8'd241;
    sbox_5[44] = 8'd113;
    sbox_5[45] = 8'd216;
    sbox_5[46] = 8'd49;
    sbox_5[47] = 8'd21;
    sbox_5[48] = 8'd4;
    sbox_5[49] = 8'd199;
    sbox_5[50] = 8'd35;
    sbox_5[51] = 8'd195;
    sbox_5[52] = 8'd24;
    sbox_5[53] = 8'd150;
    sbox_5[54] = 8'd5;
    sbox_5[55] = 8'd154;
    sbox_5[56] = 8'd7;
    sbox_5[57] = 8'd18;
    sbox_5[58] = 8'd128;
    sbox_5[59] = 8'd226;
    sbox_5[60] = 8'd235;
    sbox_5[61] = 8'd39;
    sbox_5[62] = 8'd178;
    sbox_5[63] = 8'd117;
    sbox_5[64] = 8'd9;
    sbox_5[65] = 8'd131;
    sbox_5[66] = 8'd44;
    sbox_5[67] = 8'd26;
    sbox_5[68] = 8'd27;
    sbox_5[69] = 8'd110;
    sbox_5[70] = 8'd90;
    sbox_5[71] = 8'd160;
    sbox_5[72] = 8'd82;
    sbox_5[73] = 8'd59;
    sbox_5[74] = 8'd214;
    sbox_5[75] = 8'd179;
    sbox_5[76] = 8'd41;
    sbox_5[77] = 8'd227;
    sbox_5[78] = 8'd47;
    sbox_5[79] = 8'd132;
    sbox_5[80] = 8'd83;
    sbox_5[81] = 8'd209;
    sbox_5[82] = 8'd0;
    sbox_5[83] = 8'd237;
    sbox_5[84] = 8'd32;
    sbox_5[85] = 8'd252;
    sbox_5[86] = 8'd177;
    sbox_5[87] = 8'd91;
    sbox_5[88] = 8'd106;
    sbox_5[89] = 8'd203;
    sbox_5[90] = 8'd190;
    sbox_5[91] = 8'd57;
    sbox_5[92] = 8'd74;
    sbox_5[93] = 8'd76;
    sbox_5[94] = 8'd88;
    sbox_5[95] = 8'd207;
    sbox_5[96] = 8'd208;
    sbox_5[97] = 8'd239;
    sbox_5[98] = 8'd170;
    sbox_5[99] = 8'd251;
    sbox_5[100] = 8'd67;
    sbox_5[101] = 8'd77;
    sbox_5[102] = 8'd51;
    sbox_5[103] = 8'd133;
    sbox_5[104] = 8'd69;
    sbox_5[105] = 8'd249;
    sbox_5[106] = 8'd2;
    sbox_5[107] = 8'd127;
    sbox_5[108] = 8'd80;
    sbox_5[109] = 8'd60;
    sbox_5[110] = 8'd159;
    sbox_5[111] = 8'd168;
    sbox_5[112] = 8'd81;
    sbox_5[113] = 8'd163;
    sbox_5[114] = 8'd64;
    sbox_5[115] = 8'd143;
    sbox_5[116] = 8'd146;
    sbox_5[117] = 8'd157;
    sbox_5[118] = 8'd56;
    sbox_5[119] = 8'd245;
    sbox_5[120] = 8'd188;
    sbox_5[121] = 8'd182;
    sbox_5[122] = 8'd218;
    sbox_5[123] = 8'd33;
    sbox_5[124] = 8'd16;
    sbox_5[125] = 8'd255;
    sbox_5[126] = 8'd243;
    sbox_5[127] = 8'd210;
    sbox_5[128] = 8'd205;
    sbox_5[129] = 8'd12;
    sbox_5[130] = 8'd19;
    sbox_5[131] = 8'd236;
    sbox_5[132] = 8'd95;
    sbox_5[133] = 8'd151;
    sbox_5[134] = 8'd68;
    sbox_5[135] = 8'd23;
    sbox_5[136] = 8'd196;
    sbox_5[137] = 8'd167;
    sbox_5[138] = 8'd126;
    sbox_5[139] = 8'd61;
    sbox_5[140] = 8'd100;
    sbox_5[141] = 8'd93;
    sbox_5[142] = 8'd25;
    sbox_5[143] = 8'd115;
    sbox_5[144] = 8'd96;
    sbox_5[145] = 8'd129;
    sbox_5[146] = 8'd79;
    sbox_5[147] = 8'd220;
    sbox_5[148] = 8'd34;
    sbox_5[149] = 8'd42;
    sbox_5[150] = 8'd144;
    sbox_5[151] = 8'd136;
    sbox_5[152] = 8'd70;
    sbox_5[153] = 8'd238;
    sbox_5[154] = 8'd184;
    sbox_5[155] = 8'd20;
    sbox_5[156] = 8'd222;
    sbox_5[157] = 8'd94;
    sbox_5[158] = 8'd11;
    sbox_5[159] = 8'd219;
    sbox_5[160] = 8'd224;
    sbox_5[161] = 8'd50;
    sbox_5[162] = 8'd58;
    sbox_5[163] = 8'd10;
    sbox_5[164] = 8'd73;
    sbox_5[165] = 8'd6;
    sbox_5[166] = 8'd36;
    sbox_5[167] = 8'd92;
    sbox_5[168] = 8'd194;
    sbox_5[169] = 8'd211;
    sbox_5[170] = 8'd172;
    sbox_5[171] = 8'd98;
    sbox_5[172] = 8'd145;
    sbox_5[173] = 8'd149;
    sbox_5[174] = 8'd228;
    sbox_5[175] = 8'd121;
    sbox_5[176] = 8'd231;
    sbox_5[177] = 8'd200;
    sbox_5[178] = 8'd55;
    sbox_5[179] = 8'd109;
    sbox_5[180] = 8'd141;
    sbox_5[181] = 8'd213;
    sbox_5[182] = 8'd78;
    sbox_5[183] = 8'd169;
    sbox_5[184] = 8'd108;
    sbox_5[185] = 8'd86;
    sbox_5[186] = 8'd244;
    sbox_5[187] = 8'd234;
    sbox_5[188] = 8'd101;
    sbox_5[189] = 8'd122;
    sbox_5[190] = 8'd174;
    sbox_5[191] = 8'd8;
    sbox_5[192] = 8'd186;
    sbox_5[193] = 8'd120;
    sbox_5[194] = 8'd37;
    sbox_5[195] = 8'd46;
    sbox_5[196] = 8'd28;
    sbox_5[197] = 8'd166;
    sbox_5[198] = 8'd180;
    sbox_5[199] = 8'd198;
    sbox_5[200] = 8'd232;
    sbox_5[201] = 8'd221;
    sbox_5[202] = 8'd116;
    sbox_5[203] = 8'd31;
    sbox_5[204] = 8'd75;
    sbox_5[205] = 8'd189;
    sbox_5[206] = 8'd139;
    sbox_5[207] = 8'd138;
    sbox_5[208] = 8'd112;
    sbox_5[209] = 8'd62;
    sbox_5[210] = 8'd181;
    sbox_5[211] = 8'd102;
    sbox_5[212] = 8'd72;
    sbox_5[213] = 8'd3;
    sbox_5[214] = 8'd246;
    sbox_5[215] = 8'd14;
    sbox_5[216] = 8'd97;
    sbox_5[217] = 8'd53;
    sbox_5[218] = 8'd87;
    sbox_5[219] = 8'd185;
    sbox_5[220] = 8'd134;
    sbox_5[221] = 8'd193;
    sbox_5[222] = 8'd29;
    sbox_5[223] = 8'd158;
    sbox_5[224] = 8'd225;
    sbox_5[225] = 8'd248;
    sbox_5[226] = 8'd152;
    sbox_5[227] = 8'd17;
    sbox_5[228] = 8'd105;
    sbox_5[229] = 8'd217;
    sbox_5[230] = 8'd142;
    sbox_5[231] = 8'd148;
    sbox_5[232] = 8'd155;
    sbox_5[233] = 8'd30;
    sbox_5[234] = 8'd135;
    sbox_5[235] = 8'd233;
    sbox_5[236] = 8'd206;
    sbox_5[237] = 8'd85;
    sbox_5[238] = 8'd40;
    sbox_5[239] = 8'd223;
    sbox_5[240] = 8'd140;
    sbox_5[241] = 8'd161;
    sbox_5[242] = 8'd137;
    sbox_5[243] = 8'd13;
    sbox_5[244] = 8'd191;
    sbox_5[245] = 8'd230;
    sbox_5[246] = 8'd66;
    sbox_5[247] = 8'd104;
    sbox_5[248] = 8'd65;
    sbox_5[249] = 8'd153;
    sbox_5[250] = 8'd45;
    sbox_5[251] = 8'd15;
    sbox_5[252] = 8'd176;
    sbox_5[253] = 8'd84;
    sbox_5[254] = 8'd187;
    sbox_5[255] = 8'd22;
    sbox_6[0] = 8'd99;
    sbox_6[1] = 8'd124;
    sbox_6[2] = 8'd119;
    sbox_6[3] = 8'd123;
    sbox_6[4] = 8'd242;
    sbox_6[5] = 8'd107;
    sbox_6[6] = 8'd111;
    sbox_6[7] = 8'd197;
    sbox_6[8] = 8'd48;
    sbox_6[9] = 8'd1;
    sbox_6[10] = 8'd103;
    sbox_6[11] = 8'd43;
    sbox_6[12] = 8'd254;
    sbox_6[13] = 8'd215;
    sbox_6[14] = 8'd171;
    sbox_6[15] = 8'd118;
    sbox_6[16] = 8'd202;
    sbox_6[17] = 8'd130;
    sbox_6[18] = 8'd201;
    sbox_6[19] = 8'd125;
    sbox_6[20] = 8'd250;
    sbox_6[21] = 8'd89;
    sbox_6[22] = 8'd71;
    sbox_6[23] = 8'd240;
    sbox_6[24] = 8'd173;
    sbox_6[25] = 8'd212;
    sbox_6[26] = 8'd162;
    sbox_6[27] = 8'd175;
    sbox_6[28] = 8'd156;
    sbox_6[29] = 8'd164;
    sbox_6[30] = 8'd114;
    sbox_6[31] = 8'd192;
    sbox_6[32] = 8'd183;
    sbox_6[33] = 8'd253;
    sbox_6[34] = 8'd147;
    sbox_6[35] = 8'd38;
    sbox_6[36] = 8'd54;
    sbox_6[37] = 8'd63;
    sbox_6[38] = 8'd247;
    sbox_6[39] = 8'd204;
    sbox_6[40] = 8'd52;
    sbox_6[41] = 8'd165;
    sbox_6[42] = 8'd229;
    sbox_6[43] = 8'd241;
    sbox_6[44] = 8'd113;
    sbox_6[45] = 8'd216;
    sbox_6[46] = 8'd49;
    sbox_6[47] = 8'd21;
    sbox_6[48] = 8'd4;
    sbox_6[49] = 8'd199;
    sbox_6[50] = 8'd35;
    sbox_6[51] = 8'd195;
    sbox_6[52] = 8'd24;
    sbox_6[53] = 8'd150;
    sbox_6[54] = 8'd5;
    sbox_6[55] = 8'd154;
    sbox_6[56] = 8'd7;
    sbox_6[57] = 8'd18;
    sbox_6[58] = 8'd128;
    sbox_6[59] = 8'd226;
    sbox_6[60] = 8'd235;
    sbox_6[61] = 8'd39;
    sbox_6[62] = 8'd178;
    sbox_6[63] = 8'd117;
    sbox_6[64] = 8'd9;
    sbox_6[65] = 8'd131;
    sbox_6[66] = 8'd44;
    sbox_6[67] = 8'd26;
    sbox_6[68] = 8'd27;
    sbox_6[69] = 8'd110;
    sbox_6[70] = 8'd90;
    sbox_6[71] = 8'd160;
    sbox_6[72] = 8'd82;
    sbox_6[73] = 8'd59;
    sbox_6[74] = 8'd214;
    sbox_6[75] = 8'd179;
    sbox_6[76] = 8'd41;
    sbox_6[77] = 8'd227;
    sbox_6[78] = 8'd47;
    sbox_6[79] = 8'd132;
    sbox_6[80] = 8'd83;
    sbox_6[81] = 8'd209;
    sbox_6[82] = 8'd0;
    sbox_6[83] = 8'd237;
    sbox_6[84] = 8'd32;
    sbox_6[85] = 8'd252;
    sbox_6[86] = 8'd177;
    sbox_6[87] = 8'd91;
    sbox_6[88] = 8'd106;
    sbox_6[89] = 8'd203;
    sbox_6[90] = 8'd190;
    sbox_6[91] = 8'd57;
    sbox_6[92] = 8'd74;
    sbox_6[93] = 8'd76;
    sbox_6[94] = 8'd88;
    sbox_6[95] = 8'd207;
    sbox_6[96] = 8'd208;
    sbox_6[97] = 8'd239;
    sbox_6[98] = 8'd170;
    sbox_6[99] = 8'd251;
    sbox_6[100] = 8'd67;
    sbox_6[101] = 8'd77;
    sbox_6[102] = 8'd51;
    sbox_6[103] = 8'd133;
    sbox_6[104] = 8'd69;
    sbox_6[105] = 8'd249;
    sbox_6[106] = 8'd2;
    sbox_6[107] = 8'd127;
    sbox_6[108] = 8'd80;
    sbox_6[109] = 8'd60;
    sbox_6[110] = 8'd159;
    sbox_6[111] = 8'd168;
    sbox_6[112] = 8'd81;
    sbox_6[113] = 8'd163;
    sbox_6[114] = 8'd64;
    sbox_6[115] = 8'd143;
    sbox_6[116] = 8'd146;
    sbox_6[117] = 8'd157;
    sbox_6[118] = 8'd56;
    sbox_6[119] = 8'd245;
    sbox_6[120] = 8'd188;
    sbox_6[121] = 8'd182;
    sbox_6[122] = 8'd218;
    sbox_6[123] = 8'd33;
    sbox_6[124] = 8'd16;
    sbox_6[125] = 8'd255;
    sbox_6[126] = 8'd243;
    sbox_6[127] = 8'd210;
    sbox_6[128] = 8'd205;
    sbox_6[129] = 8'd12;
    sbox_6[130] = 8'd19;
    sbox_6[131] = 8'd236;
    sbox_6[132] = 8'd95;
    sbox_6[133] = 8'd151;
    sbox_6[134] = 8'd68;
    sbox_6[135] = 8'd23;
    sbox_6[136] = 8'd196;
    sbox_6[137] = 8'd167;
    sbox_6[138] = 8'd126;
    sbox_6[139] = 8'd61;
    sbox_6[140] = 8'd100;
    sbox_6[141] = 8'd93;
    sbox_6[142] = 8'd25;
    sbox_6[143] = 8'd115;
    sbox_6[144] = 8'd96;
    sbox_6[145] = 8'd129;
    sbox_6[146] = 8'd79;
    sbox_6[147] = 8'd220;
    sbox_6[148] = 8'd34;
    sbox_6[149] = 8'd42;
    sbox_6[150] = 8'd144;
    sbox_6[151] = 8'd136;
    sbox_6[152] = 8'd70;
    sbox_6[153] = 8'd238;
    sbox_6[154] = 8'd184;
    sbox_6[155] = 8'd20;
    sbox_6[156] = 8'd222;
    sbox_6[157] = 8'd94;
    sbox_6[158] = 8'd11;
    sbox_6[159] = 8'd219;
    sbox_6[160] = 8'd224;
    sbox_6[161] = 8'd50;
    sbox_6[162] = 8'd58;
    sbox_6[163] = 8'd10;
    sbox_6[164] = 8'd73;
    sbox_6[165] = 8'd6;
    sbox_6[166] = 8'd36;
    sbox_6[167] = 8'd92;
    sbox_6[168] = 8'd194;
    sbox_6[169] = 8'd211;
    sbox_6[170] = 8'd172;
    sbox_6[171] = 8'd98;
    sbox_6[172] = 8'd145;
    sbox_6[173] = 8'd149;
    sbox_6[174] = 8'd228;
    sbox_6[175] = 8'd121;
    sbox_6[176] = 8'd231;
    sbox_6[177] = 8'd200;
    sbox_6[178] = 8'd55;
    sbox_6[179] = 8'd109;
    sbox_6[180] = 8'd141;
    sbox_6[181] = 8'd213;
    sbox_6[182] = 8'd78;
    sbox_6[183] = 8'd169;
    sbox_6[184] = 8'd108;
    sbox_6[185] = 8'd86;
    sbox_6[186] = 8'd244;
    sbox_6[187] = 8'd234;
    sbox_6[188] = 8'd101;
    sbox_6[189] = 8'd122;
    sbox_6[190] = 8'd174;
    sbox_6[191] = 8'd8;
    sbox_6[192] = 8'd186;
    sbox_6[193] = 8'd120;
    sbox_6[194] = 8'd37;
    sbox_6[195] = 8'd46;
    sbox_6[196] = 8'd28;
    sbox_6[197] = 8'd166;
    sbox_6[198] = 8'd180;
    sbox_6[199] = 8'd198;
    sbox_6[200] = 8'd232;
    sbox_6[201] = 8'd221;
    sbox_6[202] = 8'd116;
    sbox_6[203] = 8'd31;
    sbox_6[204] = 8'd75;
    sbox_6[205] = 8'd189;
    sbox_6[206] = 8'd139;
    sbox_6[207] = 8'd138;
    sbox_6[208] = 8'd112;
    sbox_6[209] = 8'd62;
    sbox_6[210] = 8'd181;
    sbox_6[211] = 8'd102;
    sbox_6[212] = 8'd72;
    sbox_6[213] = 8'd3;
    sbox_6[214] = 8'd246;
    sbox_6[215] = 8'd14;
    sbox_6[216] = 8'd97;
    sbox_6[217] = 8'd53;
    sbox_6[218] = 8'd87;
    sbox_6[219] = 8'd185;
    sbox_6[220] = 8'd134;
    sbox_6[221] = 8'd193;
    sbox_6[222] = 8'd29;
    sbox_6[223] = 8'd158;
    sbox_6[224] = 8'd225;
    sbox_6[225] = 8'd248;
    sbox_6[226] = 8'd152;
    sbox_6[227] = 8'd17;
    sbox_6[228] = 8'd105;
    sbox_6[229] = 8'd217;
    sbox_6[230] = 8'd142;
    sbox_6[231] = 8'd148;
    sbox_6[232] = 8'd155;
    sbox_6[233] = 8'd30;
    sbox_6[234] = 8'd135;
    sbox_6[235] = 8'd233;
    sbox_6[236] = 8'd206;
    sbox_6[237] = 8'd85;
    sbox_6[238] = 8'd40;
    sbox_6[239] = 8'd223;
    sbox_6[240] = 8'd140;
    sbox_6[241] = 8'd161;
    sbox_6[242] = 8'd137;
    sbox_6[243] = 8'd13;
    sbox_6[244] = 8'd191;
    sbox_6[245] = 8'd230;
    sbox_6[246] = 8'd66;
    sbox_6[247] = 8'd104;
    sbox_6[248] = 8'd65;
    sbox_6[249] = 8'd153;
    sbox_6[250] = 8'd45;
    sbox_6[251] = 8'd15;
    sbox_6[252] = 8'd176;
    sbox_6[253] = 8'd84;
    sbox_6[254] = 8'd187;
    sbox_6[255] = 8'd22;
    sbox_7[0] = 8'd99;
    sbox_7[1] = 8'd124;
    sbox_7[2] = 8'd119;
    sbox_7[3] = 8'd123;
    sbox_7[4] = 8'd242;
    sbox_7[5] = 8'd107;
    sbox_7[6] = 8'd111;
    sbox_7[7] = 8'd197;
    sbox_7[8] = 8'd48;
    sbox_7[9] = 8'd1;
    sbox_7[10] = 8'd103;
    sbox_7[11] = 8'd43;
    sbox_7[12] = 8'd254;
    sbox_7[13] = 8'd215;
    sbox_7[14] = 8'd171;
    sbox_7[15] = 8'd118;
    sbox_7[16] = 8'd202;
    sbox_7[17] = 8'd130;
    sbox_7[18] = 8'd201;
    sbox_7[19] = 8'd125;
    sbox_7[20] = 8'd250;
    sbox_7[21] = 8'd89;
    sbox_7[22] = 8'd71;
    sbox_7[23] = 8'd240;
    sbox_7[24] = 8'd173;
    sbox_7[25] = 8'd212;
    sbox_7[26] = 8'd162;
    sbox_7[27] = 8'd175;
    sbox_7[28] = 8'd156;
    sbox_7[29] = 8'd164;
    sbox_7[30] = 8'd114;
    sbox_7[31] = 8'd192;
    sbox_7[32] = 8'd183;
    sbox_7[33] = 8'd253;
    sbox_7[34] = 8'd147;
    sbox_7[35] = 8'd38;
    sbox_7[36] = 8'd54;
    sbox_7[37] = 8'd63;
    sbox_7[38] = 8'd247;
    sbox_7[39] = 8'd204;
    sbox_7[40] = 8'd52;
    sbox_7[41] = 8'd165;
    sbox_7[42] = 8'd229;
    sbox_7[43] = 8'd241;
    sbox_7[44] = 8'd113;
    sbox_7[45] = 8'd216;
    sbox_7[46] = 8'd49;
    sbox_7[47] = 8'd21;
    sbox_7[48] = 8'd4;
    sbox_7[49] = 8'd199;
    sbox_7[50] = 8'd35;
    sbox_7[51] = 8'd195;
    sbox_7[52] = 8'd24;
    sbox_7[53] = 8'd150;
    sbox_7[54] = 8'd5;
    sbox_7[55] = 8'd154;
    sbox_7[56] = 8'd7;
    sbox_7[57] = 8'd18;
    sbox_7[58] = 8'd128;
    sbox_7[59] = 8'd226;
    sbox_7[60] = 8'd235;
    sbox_7[61] = 8'd39;
    sbox_7[62] = 8'd178;
    sbox_7[63] = 8'd117;
    sbox_7[64] = 8'd9;
    sbox_7[65] = 8'd131;
    sbox_7[66] = 8'd44;
    sbox_7[67] = 8'd26;
    sbox_7[68] = 8'd27;
    sbox_7[69] = 8'd110;
    sbox_7[70] = 8'd90;
    sbox_7[71] = 8'd160;
    sbox_7[72] = 8'd82;
    sbox_7[73] = 8'd59;
    sbox_7[74] = 8'd214;
    sbox_7[75] = 8'd179;
    sbox_7[76] = 8'd41;
    sbox_7[77] = 8'd227;
    sbox_7[78] = 8'd47;
    sbox_7[79] = 8'd132;
    sbox_7[80] = 8'd83;
    sbox_7[81] = 8'd209;
    sbox_7[82] = 8'd0;
    sbox_7[83] = 8'd237;
    sbox_7[84] = 8'd32;
    sbox_7[85] = 8'd252;
    sbox_7[86] = 8'd177;
    sbox_7[87] = 8'd91;
    sbox_7[88] = 8'd106;
    sbox_7[89] = 8'd203;
    sbox_7[90] = 8'd190;
    sbox_7[91] = 8'd57;
    sbox_7[92] = 8'd74;
    sbox_7[93] = 8'd76;
    sbox_7[94] = 8'd88;
    sbox_7[95] = 8'd207;
    sbox_7[96] = 8'd208;
    sbox_7[97] = 8'd239;
    sbox_7[98] = 8'd170;
    sbox_7[99] = 8'd251;
    sbox_7[100] = 8'd67;
    sbox_7[101] = 8'd77;
    sbox_7[102] = 8'd51;
    sbox_7[103] = 8'd133;
    sbox_7[104] = 8'd69;
    sbox_7[105] = 8'd249;
    sbox_7[106] = 8'd2;
    sbox_7[107] = 8'd127;
    sbox_7[108] = 8'd80;
    sbox_7[109] = 8'd60;
    sbox_7[110] = 8'd159;
    sbox_7[111] = 8'd168;
    sbox_7[112] = 8'd81;
    sbox_7[113] = 8'd163;
    sbox_7[114] = 8'd64;
    sbox_7[115] = 8'd143;
    sbox_7[116] = 8'd146;
    sbox_7[117] = 8'd157;
    sbox_7[118] = 8'd56;
    sbox_7[119] = 8'd245;
    sbox_7[120] = 8'd188;
    sbox_7[121] = 8'd182;
    sbox_7[122] = 8'd218;
    sbox_7[123] = 8'd33;
    sbox_7[124] = 8'd16;
    sbox_7[125] = 8'd255;
    sbox_7[126] = 8'd243;
    sbox_7[127] = 8'd210;
    sbox_7[128] = 8'd205;
    sbox_7[129] = 8'd12;
    sbox_7[130] = 8'd19;
    sbox_7[131] = 8'd236;
    sbox_7[132] = 8'd95;
    sbox_7[133] = 8'd151;
    sbox_7[134] = 8'd68;
    sbox_7[135] = 8'd23;
    sbox_7[136] = 8'd196;
    sbox_7[137] = 8'd167;
    sbox_7[138] = 8'd126;
    sbox_7[139] = 8'd61;
    sbox_7[140] = 8'd100;
    sbox_7[141] = 8'd93;
    sbox_7[142] = 8'd25;
    sbox_7[143] = 8'd115;
    sbox_7[144] = 8'd96;
    sbox_7[145] = 8'd129;
    sbox_7[146] = 8'd79;
    sbox_7[147] = 8'd220;
    sbox_7[148] = 8'd34;
    sbox_7[149] = 8'd42;
    sbox_7[150] = 8'd144;
    sbox_7[151] = 8'd136;
    sbox_7[152] = 8'd70;
    sbox_7[153] = 8'd238;
    sbox_7[154] = 8'd184;
    sbox_7[155] = 8'd20;
    sbox_7[156] = 8'd222;
    sbox_7[157] = 8'd94;
    sbox_7[158] = 8'd11;
    sbox_7[159] = 8'd219;
    sbox_7[160] = 8'd224;
    sbox_7[161] = 8'd50;
    sbox_7[162] = 8'd58;
    sbox_7[163] = 8'd10;
    sbox_7[164] = 8'd73;
    sbox_7[165] = 8'd6;
    sbox_7[166] = 8'd36;
    sbox_7[167] = 8'd92;
    sbox_7[168] = 8'd194;
    sbox_7[169] = 8'd211;
    sbox_7[170] = 8'd172;
    sbox_7[171] = 8'd98;
    sbox_7[172] = 8'd145;
    sbox_7[173] = 8'd149;
    sbox_7[174] = 8'd228;
    sbox_7[175] = 8'd121;
    sbox_7[176] = 8'd231;
    sbox_7[177] = 8'd200;
    sbox_7[178] = 8'd55;
    sbox_7[179] = 8'd109;
    sbox_7[180] = 8'd141;
    sbox_7[181] = 8'd213;
    sbox_7[182] = 8'd78;
    sbox_7[183] = 8'd169;
    sbox_7[184] = 8'd108;
    sbox_7[185] = 8'd86;
    sbox_7[186] = 8'd244;
    sbox_7[187] = 8'd234;
    sbox_7[188] = 8'd101;
    sbox_7[189] = 8'd122;
    sbox_7[190] = 8'd174;
    sbox_7[191] = 8'd8;
    sbox_7[192] = 8'd186;
    sbox_7[193] = 8'd120;
    sbox_7[194] = 8'd37;
    sbox_7[195] = 8'd46;
    sbox_7[196] = 8'd28;
    sbox_7[197] = 8'd166;
    sbox_7[198] = 8'd180;
    sbox_7[199] = 8'd198;
    sbox_7[200] = 8'd232;
    sbox_7[201] = 8'd221;
    sbox_7[202] = 8'd116;
    sbox_7[203] = 8'd31;
    sbox_7[204] = 8'd75;
    sbox_7[205] = 8'd189;
    sbox_7[206] = 8'd139;
    sbox_7[207] = 8'd138;
    sbox_7[208] = 8'd112;
    sbox_7[209] = 8'd62;
    sbox_7[210] = 8'd181;
    sbox_7[211] = 8'd102;
    sbox_7[212] = 8'd72;
    sbox_7[213] = 8'd3;
    sbox_7[214] = 8'd246;
    sbox_7[215] = 8'd14;
    sbox_7[216] = 8'd97;
    sbox_7[217] = 8'd53;
    sbox_7[218] = 8'd87;
    sbox_7[219] = 8'd185;
    sbox_7[220] = 8'd134;
    sbox_7[221] = 8'd193;
    sbox_7[222] = 8'd29;
    sbox_7[223] = 8'd158;
    sbox_7[224] = 8'd225;
    sbox_7[225] = 8'd248;
    sbox_7[226] = 8'd152;
    sbox_7[227] = 8'd17;
    sbox_7[228] = 8'd105;
    sbox_7[229] = 8'd217;
    sbox_7[230] = 8'd142;
    sbox_7[231] = 8'd148;
    sbox_7[232] = 8'd155;
    sbox_7[233] = 8'd30;
    sbox_7[234] = 8'd135;
    sbox_7[235] = 8'd233;
    sbox_7[236] = 8'd206;
    sbox_7[237] = 8'd85;
    sbox_7[238] = 8'd40;
    sbox_7[239] = 8'd223;
    sbox_7[240] = 8'd140;
    sbox_7[241] = 8'd161;
    sbox_7[242] = 8'd137;
    sbox_7[243] = 8'd13;
    sbox_7[244] = 8'd191;
    sbox_7[245] = 8'd230;
    sbox_7[246] = 8'd66;
    sbox_7[247] = 8'd104;
    sbox_7[248] = 8'd65;
    sbox_7[249] = 8'd153;
    sbox_7[250] = 8'd45;
    sbox_7[251] = 8'd15;
    sbox_7[252] = 8'd176;
    sbox_7[253] = 8'd84;
    sbox_7[254] = 8'd187;
    sbox_7[255] = 8'd22;
    sbox_8[0] = 8'd99;
    sbox_8[1] = 8'd124;
    sbox_8[2] = 8'd119;
    sbox_8[3] = 8'd123;
    sbox_8[4] = 8'd242;
    sbox_8[5] = 8'd107;
    sbox_8[6] = 8'd111;
    sbox_8[7] = 8'd197;
    sbox_8[8] = 8'd48;
    sbox_8[9] = 8'd1;
    sbox_8[10] = 8'd103;
    sbox_8[11] = 8'd43;
    sbox_8[12] = 8'd254;
    sbox_8[13] = 8'd215;
    sbox_8[14] = 8'd171;
    sbox_8[15] = 8'd118;
    sbox_8[16] = 8'd202;
    sbox_8[17] = 8'd130;
    sbox_8[18] = 8'd201;
    sbox_8[19] = 8'd125;
    sbox_8[20] = 8'd250;
    sbox_8[21] = 8'd89;
    sbox_8[22] = 8'd71;
    sbox_8[23] = 8'd240;
    sbox_8[24] = 8'd173;
    sbox_8[25] = 8'd212;
    sbox_8[26] = 8'd162;
    sbox_8[27] = 8'd175;
    sbox_8[28] = 8'd156;
    sbox_8[29] = 8'd164;
    sbox_8[30] = 8'd114;
    sbox_8[31] = 8'd192;
    sbox_8[32] = 8'd183;
    sbox_8[33] = 8'd253;
    sbox_8[34] = 8'd147;
    sbox_8[35] = 8'd38;
    sbox_8[36] = 8'd54;
    sbox_8[37] = 8'd63;
    sbox_8[38] = 8'd247;
    sbox_8[39] = 8'd204;
    sbox_8[40] = 8'd52;
    sbox_8[41] = 8'd165;
    sbox_8[42] = 8'd229;
    sbox_8[43] = 8'd241;
    sbox_8[44] = 8'd113;
    sbox_8[45] = 8'd216;
    sbox_8[46] = 8'd49;
    sbox_8[47] = 8'd21;
    sbox_8[48] = 8'd4;
    sbox_8[49] = 8'd199;
    sbox_8[50] = 8'd35;
    sbox_8[51] = 8'd195;
    sbox_8[52] = 8'd24;
    sbox_8[53] = 8'd150;
    sbox_8[54] = 8'd5;
    sbox_8[55] = 8'd154;
    sbox_8[56] = 8'd7;
    sbox_8[57] = 8'd18;
    sbox_8[58] = 8'd128;
    sbox_8[59] = 8'd226;
    sbox_8[60] = 8'd235;
    sbox_8[61] = 8'd39;
    sbox_8[62] = 8'd178;
    sbox_8[63] = 8'd117;
    sbox_8[64] = 8'd9;
    sbox_8[65] = 8'd131;
    sbox_8[66] = 8'd44;
    sbox_8[67] = 8'd26;
    sbox_8[68] = 8'd27;
    sbox_8[69] = 8'd110;
    sbox_8[70] = 8'd90;
    sbox_8[71] = 8'd160;
    sbox_8[72] = 8'd82;
    sbox_8[73] = 8'd59;
    sbox_8[74] = 8'd214;
    sbox_8[75] = 8'd179;
    sbox_8[76] = 8'd41;
    sbox_8[77] = 8'd227;
    sbox_8[78] = 8'd47;
    sbox_8[79] = 8'd132;
    sbox_8[80] = 8'd83;
    sbox_8[81] = 8'd209;
    sbox_8[82] = 8'd0;
    sbox_8[83] = 8'd237;
    sbox_8[84] = 8'd32;
    sbox_8[85] = 8'd252;
    sbox_8[86] = 8'd177;
    sbox_8[87] = 8'd91;
    sbox_8[88] = 8'd106;
    sbox_8[89] = 8'd203;
    sbox_8[90] = 8'd190;
    sbox_8[91] = 8'd57;
    sbox_8[92] = 8'd74;
    sbox_8[93] = 8'd76;
    sbox_8[94] = 8'd88;
    sbox_8[95] = 8'd207;
    sbox_8[96] = 8'd208;
    sbox_8[97] = 8'd239;
    sbox_8[98] = 8'd170;
    sbox_8[99] = 8'd251;
    sbox_8[100] = 8'd67;
    sbox_8[101] = 8'd77;
    sbox_8[102] = 8'd51;
    sbox_8[103] = 8'd133;
    sbox_8[104] = 8'd69;
    sbox_8[105] = 8'd249;
    sbox_8[106] = 8'd2;
    sbox_8[107] = 8'd127;
    sbox_8[108] = 8'd80;
    sbox_8[109] = 8'd60;
    sbox_8[110] = 8'd159;
    sbox_8[111] = 8'd168;
    sbox_8[112] = 8'd81;
    sbox_8[113] = 8'd163;
    sbox_8[114] = 8'd64;
    sbox_8[115] = 8'd143;
    sbox_8[116] = 8'd146;
    sbox_8[117] = 8'd157;
    sbox_8[118] = 8'd56;
    sbox_8[119] = 8'd245;
    sbox_8[120] = 8'd188;
    sbox_8[121] = 8'd182;
    sbox_8[122] = 8'd218;
    sbox_8[123] = 8'd33;
    sbox_8[124] = 8'd16;
    sbox_8[125] = 8'd255;
    sbox_8[126] = 8'd243;
    sbox_8[127] = 8'd210;
    sbox_8[128] = 8'd205;
    sbox_8[129] = 8'd12;
    sbox_8[130] = 8'd19;
    sbox_8[131] = 8'd236;
    sbox_8[132] = 8'd95;
    sbox_8[133] = 8'd151;
    sbox_8[134] = 8'd68;
    sbox_8[135] = 8'd23;
    sbox_8[136] = 8'd196;
    sbox_8[137] = 8'd167;
    sbox_8[138] = 8'd126;
    sbox_8[139] = 8'd61;
    sbox_8[140] = 8'd100;
    sbox_8[141] = 8'd93;
    sbox_8[142] = 8'd25;
    sbox_8[143] = 8'd115;
    sbox_8[144] = 8'd96;
    sbox_8[145] = 8'd129;
    sbox_8[146] = 8'd79;
    sbox_8[147] = 8'd220;
    sbox_8[148] = 8'd34;
    sbox_8[149] = 8'd42;
    sbox_8[150] = 8'd144;
    sbox_8[151] = 8'd136;
    sbox_8[152] = 8'd70;
    sbox_8[153] = 8'd238;
    sbox_8[154] = 8'd184;
    sbox_8[155] = 8'd20;
    sbox_8[156] = 8'd222;
    sbox_8[157] = 8'd94;
    sbox_8[158] = 8'd11;
    sbox_8[159] = 8'd219;
    sbox_8[160] = 8'd224;
    sbox_8[161] = 8'd50;
    sbox_8[162] = 8'd58;
    sbox_8[163] = 8'd10;
    sbox_8[164] = 8'd73;
    sbox_8[165] = 8'd6;
    sbox_8[166] = 8'd36;
    sbox_8[167] = 8'd92;
    sbox_8[168] = 8'd194;
    sbox_8[169] = 8'd211;
    sbox_8[170] = 8'd172;
    sbox_8[171] = 8'd98;
    sbox_8[172] = 8'd145;
    sbox_8[173] = 8'd149;
    sbox_8[174] = 8'd228;
    sbox_8[175] = 8'd121;
    sbox_8[176] = 8'd231;
    sbox_8[177] = 8'd200;
    sbox_8[178] = 8'd55;
    sbox_8[179] = 8'd109;
    sbox_8[180] = 8'd141;
    sbox_8[181] = 8'd213;
    sbox_8[182] = 8'd78;
    sbox_8[183] = 8'd169;
    sbox_8[184] = 8'd108;
    sbox_8[185] = 8'd86;
    sbox_8[186] = 8'd244;
    sbox_8[187] = 8'd234;
    sbox_8[188] = 8'd101;
    sbox_8[189] = 8'd122;
    sbox_8[190] = 8'd174;
    sbox_8[191] = 8'd8;
    sbox_8[192] = 8'd186;
    sbox_8[193] = 8'd120;
    sbox_8[194] = 8'd37;
    sbox_8[195] = 8'd46;
    sbox_8[196] = 8'd28;
    sbox_8[197] = 8'd166;
    sbox_8[198] = 8'd180;
    sbox_8[199] = 8'd198;
    sbox_8[200] = 8'd232;
    sbox_8[201] = 8'd221;
    sbox_8[202] = 8'd116;
    sbox_8[203] = 8'd31;
    sbox_8[204] = 8'd75;
    sbox_8[205] = 8'd189;
    sbox_8[206] = 8'd139;
    sbox_8[207] = 8'd138;
    sbox_8[208] = 8'd112;
    sbox_8[209] = 8'd62;
    sbox_8[210] = 8'd181;
    sbox_8[211] = 8'd102;
    sbox_8[212] = 8'd72;
    sbox_8[213] = 8'd3;
    sbox_8[214] = 8'd246;
    sbox_8[215] = 8'd14;
    sbox_8[216] = 8'd97;
    sbox_8[217] = 8'd53;
    sbox_8[218] = 8'd87;
    sbox_8[219] = 8'd185;
    sbox_8[220] = 8'd134;
    sbox_8[221] = 8'd193;
    sbox_8[222] = 8'd29;
    sbox_8[223] = 8'd158;
    sbox_8[224] = 8'd225;
    sbox_8[225] = 8'd248;
    sbox_8[226] = 8'd152;
    sbox_8[227] = 8'd17;
    sbox_8[228] = 8'd105;
    sbox_8[229] = 8'd217;
    sbox_8[230] = 8'd142;
    sbox_8[231] = 8'd148;
    sbox_8[232] = 8'd155;
    sbox_8[233] = 8'd30;
    sbox_8[234] = 8'd135;
    sbox_8[235] = 8'd233;
    sbox_8[236] = 8'd206;
    sbox_8[237] = 8'd85;
    sbox_8[238] = 8'd40;
    sbox_8[239] = 8'd223;
    sbox_8[240] = 8'd140;
    sbox_8[241] = 8'd161;
    sbox_8[242] = 8'd137;
    sbox_8[243] = 8'd13;
    sbox_8[244] = 8'd191;
    sbox_8[245] = 8'd230;
    sbox_8[246] = 8'd66;
    sbox_8[247] = 8'd104;
    sbox_8[248] = 8'd65;
    sbox_8[249] = 8'd153;
    sbox_8[250] = 8'd45;
    sbox_8[251] = 8'd15;
    sbox_8[252] = 8'd176;
    sbox_8[253] = 8'd84;
    sbox_8[254] = 8'd187;
    sbox_8[255] = 8'd22;
    sbox_9[0] = 8'd99;
    sbox_9[1] = 8'd124;
    sbox_9[2] = 8'd119;
    sbox_9[3] = 8'd123;
    sbox_9[4] = 8'd242;
    sbox_9[5] = 8'd107;
    sbox_9[6] = 8'd111;
    sbox_9[7] = 8'd197;
    sbox_9[8] = 8'd48;
    sbox_9[9] = 8'd1;
    sbox_9[10] = 8'd103;
    sbox_9[11] = 8'd43;
    sbox_9[12] = 8'd254;
    sbox_9[13] = 8'd215;
    sbox_9[14] = 8'd171;
    sbox_9[15] = 8'd118;
    sbox_9[16] = 8'd202;
    sbox_9[17] = 8'd130;
    sbox_9[18] = 8'd201;
    sbox_9[19] = 8'd125;
    sbox_9[20] = 8'd250;
    sbox_9[21] = 8'd89;
    sbox_9[22] = 8'd71;
    sbox_9[23] = 8'd240;
    sbox_9[24] = 8'd173;
    sbox_9[25] = 8'd212;
    sbox_9[26] = 8'd162;
    sbox_9[27] = 8'd175;
    sbox_9[28] = 8'd156;
    sbox_9[29] = 8'd164;
    sbox_9[30] = 8'd114;
    sbox_9[31] = 8'd192;
    sbox_9[32] = 8'd183;
    sbox_9[33] = 8'd253;
    sbox_9[34] = 8'd147;
    sbox_9[35] = 8'd38;
    sbox_9[36] = 8'd54;
    sbox_9[37] = 8'd63;
    sbox_9[38] = 8'd247;
    sbox_9[39] = 8'd204;
    sbox_9[40] = 8'd52;
    sbox_9[41] = 8'd165;
    sbox_9[42] = 8'd229;
    sbox_9[43] = 8'd241;
    sbox_9[44] = 8'd113;
    sbox_9[45] = 8'd216;
    sbox_9[46] = 8'd49;
    sbox_9[47] = 8'd21;
    sbox_9[48] = 8'd4;
    sbox_9[49] = 8'd199;
    sbox_9[50] = 8'd35;
    sbox_9[51] = 8'd195;
    sbox_9[52] = 8'd24;
    sbox_9[53] = 8'd150;
    sbox_9[54] = 8'd5;
    sbox_9[55] = 8'd154;
    sbox_9[56] = 8'd7;
    sbox_9[57] = 8'd18;
    sbox_9[58] = 8'd128;
    sbox_9[59] = 8'd226;
    sbox_9[60] = 8'd235;
    sbox_9[61] = 8'd39;
    sbox_9[62] = 8'd178;
    sbox_9[63] = 8'd117;
    sbox_9[64] = 8'd9;
    sbox_9[65] = 8'd131;
    sbox_9[66] = 8'd44;
    sbox_9[67] = 8'd26;
    sbox_9[68] = 8'd27;
    sbox_9[69] = 8'd110;
    sbox_9[70] = 8'd90;
    sbox_9[71] = 8'd160;
    sbox_9[72] = 8'd82;
    sbox_9[73] = 8'd59;
    sbox_9[74] = 8'd214;
    sbox_9[75] = 8'd179;
    sbox_9[76] = 8'd41;
    sbox_9[77] = 8'd227;
    sbox_9[78] = 8'd47;
    sbox_9[79] = 8'd132;
    sbox_9[80] = 8'd83;
    sbox_9[81] = 8'd209;
    sbox_9[82] = 8'd0;
    sbox_9[83] = 8'd237;
    sbox_9[84] = 8'd32;
    sbox_9[85] = 8'd252;
    sbox_9[86] = 8'd177;
    sbox_9[87] = 8'd91;
    sbox_9[88] = 8'd106;
    sbox_9[89] = 8'd203;
    sbox_9[90] = 8'd190;
    sbox_9[91] = 8'd57;
    sbox_9[92] = 8'd74;
    sbox_9[93] = 8'd76;
    sbox_9[94] = 8'd88;
    sbox_9[95] = 8'd207;
    sbox_9[96] = 8'd208;
    sbox_9[97] = 8'd239;
    sbox_9[98] = 8'd170;
    sbox_9[99] = 8'd251;
    sbox_9[100] = 8'd67;
    sbox_9[101] = 8'd77;
    sbox_9[102] = 8'd51;
    sbox_9[103] = 8'd133;
    sbox_9[104] = 8'd69;
    sbox_9[105] = 8'd249;
    sbox_9[106] = 8'd2;
    sbox_9[107] = 8'd127;
    sbox_9[108] = 8'd80;
    sbox_9[109] = 8'd60;
    sbox_9[110] = 8'd159;
    sbox_9[111] = 8'd168;
    sbox_9[112] = 8'd81;
    sbox_9[113] = 8'd163;
    sbox_9[114] = 8'd64;
    sbox_9[115] = 8'd143;
    sbox_9[116] = 8'd146;
    sbox_9[117] = 8'd157;
    sbox_9[118] = 8'd56;
    sbox_9[119] = 8'd245;
    sbox_9[120] = 8'd188;
    sbox_9[121] = 8'd182;
    sbox_9[122] = 8'd218;
    sbox_9[123] = 8'd33;
    sbox_9[124] = 8'd16;
    sbox_9[125] = 8'd255;
    sbox_9[126] = 8'd243;
    sbox_9[127] = 8'd210;
    sbox_9[128] = 8'd205;
    sbox_9[129] = 8'd12;
    sbox_9[130] = 8'd19;
    sbox_9[131] = 8'd236;
    sbox_9[132] = 8'd95;
    sbox_9[133] = 8'd151;
    sbox_9[134] = 8'd68;
    sbox_9[135] = 8'd23;
    sbox_9[136] = 8'd196;
    sbox_9[137] = 8'd167;
    sbox_9[138] = 8'd126;
    sbox_9[139] = 8'd61;
    sbox_9[140] = 8'd100;
    sbox_9[141] = 8'd93;
    sbox_9[142] = 8'd25;
    sbox_9[143] = 8'd115;
    sbox_9[144] = 8'd96;
    sbox_9[145] = 8'd129;
    sbox_9[146] = 8'd79;
    sbox_9[147] = 8'd220;
    sbox_9[148] = 8'd34;
    sbox_9[149] = 8'd42;
    sbox_9[150] = 8'd144;
    sbox_9[151] = 8'd136;
    sbox_9[152] = 8'd70;
    sbox_9[153] = 8'd238;
    sbox_9[154] = 8'd184;
    sbox_9[155] = 8'd20;
    sbox_9[156] = 8'd222;
    sbox_9[157] = 8'd94;
    sbox_9[158] = 8'd11;
    sbox_9[159] = 8'd219;
    sbox_9[160] = 8'd224;
    sbox_9[161] = 8'd50;
    sbox_9[162] = 8'd58;
    sbox_9[163] = 8'd10;
    sbox_9[164] = 8'd73;
    sbox_9[165] = 8'd6;
    sbox_9[166] = 8'd36;
    sbox_9[167] = 8'd92;
    sbox_9[168] = 8'd194;
    sbox_9[169] = 8'd211;
    sbox_9[170] = 8'd172;
    sbox_9[171] = 8'd98;
    sbox_9[172] = 8'd145;
    sbox_9[173] = 8'd149;
    sbox_9[174] = 8'd228;
    sbox_9[175] = 8'd121;
    sbox_9[176] = 8'd231;
    sbox_9[177] = 8'd200;
    sbox_9[178] = 8'd55;
    sbox_9[179] = 8'd109;
    sbox_9[180] = 8'd141;
    sbox_9[181] = 8'd213;
    sbox_9[182] = 8'd78;
    sbox_9[183] = 8'd169;
    sbox_9[184] = 8'd108;
    sbox_9[185] = 8'd86;
    sbox_9[186] = 8'd244;
    sbox_9[187] = 8'd234;
    sbox_9[188] = 8'd101;
    sbox_9[189] = 8'd122;
    sbox_9[190] = 8'd174;
    sbox_9[191] = 8'd8;
    sbox_9[192] = 8'd186;
    sbox_9[193] = 8'd120;
    sbox_9[194] = 8'd37;
    sbox_9[195] = 8'd46;
    sbox_9[196] = 8'd28;
    sbox_9[197] = 8'd166;
    sbox_9[198] = 8'd180;
    sbox_9[199] = 8'd198;
    sbox_9[200] = 8'd232;
    sbox_9[201] = 8'd221;
    sbox_9[202] = 8'd116;
    sbox_9[203] = 8'd31;
    sbox_9[204] = 8'd75;
    sbox_9[205] = 8'd189;
    sbox_9[206] = 8'd139;
    sbox_9[207] = 8'd138;
    sbox_9[208] = 8'd112;
    sbox_9[209] = 8'd62;
    sbox_9[210] = 8'd181;
    sbox_9[211] = 8'd102;
    sbox_9[212] = 8'd72;
    sbox_9[213] = 8'd3;
    sbox_9[214] = 8'd246;
    sbox_9[215] = 8'd14;
    sbox_9[216] = 8'd97;
    sbox_9[217] = 8'd53;
    sbox_9[218] = 8'd87;
    sbox_9[219] = 8'd185;
    sbox_9[220] = 8'd134;
    sbox_9[221] = 8'd193;
    sbox_9[222] = 8'd29;
    sbox_9[223] = 8'd158;
    sbox_9[224] = 8'd225;
    sbox_9[225] = 8'd248;
    sbox_9[226] = 8'd152;
    sbox_9[227] = 8'd17;
    sbox_9[228] = 8'd105;
    sbox_9[229] = 8'd217;
    sbox_9[230] = 8'd142;
    sbox_9[231] = 8'd148;
    sbox_9[232] = 8'd155;
    sbox_9[233] = 8'd30;
    sbox_9[234] = 8'd135;
    sbox_9[235] = 8'd233;
    sbox_9[236] = 8'd206;
    sbox_9[237] = 8'd85;
    sbox_9[238] = 8'd40;
    sbox_9[239] = 8'd223;
    sbox_9[240] = 8'd140;
    sbox_9[241] = 8'd161;
    sbox_9[242] = 8'd137;
    sbox_9[243] = 8'd13;
    sbox_9[244] = 8'd191;
    sbox_9[245] = 8'd230;
    sbox_9[246] = 8'd66;
    sbox_9[247] = 8'd104;
    sbox_9[248] = 8'd65;
    sbox_9[249] = 8'd153;
    sbox_9[250] = 8'd45;
    sbox_9[251] = 8'd15;
    sbox_9[252] = 8'd176;
    sbox_9[253] = 8'd84;
    sbox_9[254] = 8'd187;
    sbox_9[255] = 8'd22;
    sbox_10[0] = 8'd99;
    sbox_10[1] = 8'd124;
    sbox_10[2] = 8'd119;
    sbox_10[3] = 8'd123;
    sbox_10[4] = 8'd242;
    sbox_10[5] = 8'd107;
    sbox_10[6] = 8'd111;
    sbox_10[7] = 8'd197;
    sbox_10[8] = 8'd48;
    sbox_10[9] = 8'd1;
    sbox_10[10] = 8'd103;
    sbox_10[11] = 8'd43;
    sbox_10[12] = 8'd254;
    sbox_10[13] = 8'd215;
    sbox_10[14] = 8'd171;
    sbox_10[15] = 8'd118;
    sbox_10[16] = 8'd202;
    sbox_10[17] = 8'd130;
    sbox_10[18] = 8'd201;
    sbox_10[19] = 8'd125;
    sbox_10[20] = 8'd250;
    sbox_10[21] = 8'd89;
    sbox_10[22] = 8'd71;
    sbox_10[23] = 8'd240;
    sbox_10[24] = 8'd173;
    sbox_10[25] = 8'd212;
    sbox_10[26] = 8'd162;
    sbox_10[27] = 8'd175;
    sbox_10[28] = 8'd156;
    sbox_10[29] = 8'd164;
    sbox_10[30] = 8'd114;
    sbox_10[31] = 8'd192;
    sbox_10[32] = 8'd183;
    sbox_10[33] = 8'd253;
    sbox_10[34] = 8'd147;
    sbox_10[35] = 8'd38;
    sbox_10[36] = 8'd54;
    sbox_10[37] = 8'd63;
    sbox_10[38] = 8'd247;
    sbox_10[39] = 8'd204;
    sbox_10[40] = 8'd52;
    sbox_10[41] = 8'd165;
    sbox_10[42] = 8'd229;
    sbox_10[43] = 8'd241;
    sbox_10[44] = 8'd113;
    sbox_10[45] = 8'd216;
    sbox_10[46] = 8'd49;
    sbox_10[47] = 8'd21;
    sbox_10[48] = 8'd4;
    sbox_10[49] = 8'd199;
    sbox_10[50] = 8'd35;
    sbox_10[51] = 8'd195;
    sbox_10[52] = 8'd24;
    sbox_10[53] = 8'd150;
    sbox_10[54] = 8'd5;
    sbox_10[55] = 8'd154;
    sbox_10[56] = 8'd7;
    sbox_10[57] = 8'd18;
    sbox_10[58] = 8'd128;
    sbox_10[59] = 8'd226;
    sbox_10[60] = 8'd235;
    sbox_10[61] = 8'd39;
    sbox_10[62] = 8'd178;
    sbox_10[63] = 8'd117;
    sbox_10[64] = 8'd9;
    sbox_10[65] = 8'd131;
    sbox_10[66] = 8'd44;
    sbox_10[67] = 8'd26;
    sbox_10[68] = 8'd27;
    sbox_10[69] = 8'd110;
    sbox_10[70] = 8'd90;
    sbox_10[71] = 8'd160;
    sbox_10[72] = 8'd82;
    sbox_10[73] = 8'd59;
    sbox_10[74] = 8'd214;
    sbox_10[75] = 8'd179;
    sbox_10[76] = 8'd41;
    sbox_10[77] = 8'd227;
    sbox_10[78] = 8'd47;
    sbox_10[79] = 8'd132;
    sbox_10[80] = 8'd83;
    sbox_10[81] = 8'd209;
    sbox_10[82] = 8'd0;
    sbox_10[83] = 8'd237;
    sbox_10[84] = 8'd32;
    sbox_10[85] = 8'd252;
    sbox_10[86] = 8'd177;
    sbox_10[87] = 8'd91;
    sbox_10[88] = 8'd106;
    sbox_10[89] = 8'd203;
    sbox_10[90] = 8'd190;
    sbox_10[91] = 8'd57;
    sbox_10[92] = 8'd74;
    sbox_10[93] = 8'd76;
    sbox_10[94] = 8'd88;
    sbox_10[95] = 8'd207;
    sbox_10[96] = 8'd208;
    sbox_10[97] = 8'd239;
    sbox_10[98] = 8'd170;
    sbox_10[99] = 8'd251;
    sbox_10[100] = 8'd67;
    sbox_10[101] = 8'd77;
    sbox_10[102] = 8'd51;
    sbox_10[103] = 8'd133;
    sbox_10[104] = 8'd69;
    sbox_10[105] = 8'd249;
    sbox_10[106] = 8'd2;
    sbox_10[107] = 8'd127;
    sbox_10[108] = 8'd80;
    sbox_10[109] = 8'd60;
    sbox_10[110] = 8'd159;
    sbox_10[111] = 8'd168;
    sbox_10[112] = 8'd81;
    sbox_10[113] = 8'd163;
    sbox_10[114] = 8'd64;
    sbox_10[115] = 8'd143;
    sbox_10[116] = 8'd146;
    sbox_10[117] = 8'd157;
    sbox_10[118] = 8'd56;
    sbox_10[119] = 8'd245;
    sbox_10[120] = 8'd188;
    sbox_10[121] = 8'd182;
    sbox_10[122] = 8'd218;
    sbox_10[123] = 8'd33;
    sbox_10[124] = 8'd16;
    sbox_10[125] = 8'd255;
    sbox_10[126] = 8'd243;
    sbox_10[127] = 8'd210;
    sbox_10[128] = 8'd205;
    sbox_10[129] = 8'd12;
    sbox_10[130] = 8'd19;
    sbox_10[131] = 8'd236;
    sbox_10[132] = 8'd95;
    sbox_10[133] = 8'd151;
    sbox_10[134] = 8'd68;
    sbox_10[135] = 8'd23;
    sbox_10[136] = 8'd196;
    sbox_10[137] = 8'd167;
    sbox_10[138] = 8'd126;
    sbox_10[139] = 8'd61;
    sbox_10[140] = 8'd100;
    sbox_10[141] = 8'd93;
    sbox_10[142] = 8'd25;
    sbox_10[143] = 8'd115;
    sbox_10[144] = 8'd96;
    sbox_10[145] = 8'd129;
    sbox_10[146] = 8'd79;
    sbox_10[147] = 8'd220;
    sbox_10[148] = 8'd34;
    sbox_10[149] = 8'd42;
    sbox_10[150] = 8'd144;
    sbox_10[151] = 8'd136;
    sbox_10[152] = 8'd70;
    sbox_10[153] = 8'd238;
    sbox_10[154] = 8'd184;
    sbox_10[155] = 8'd20;
    sbox_10[156] = 8'd222;
    sbox_10[157] = 8'd94;
    sbox_10[158] = 8'd11;
    sbox_10[159] = 8'd219;
    sbox_10[160] = 8'd224;
    sbox_10[161] = 8'd50;
    sbox_10[162] = 8'd58;
    sbox_10[163] = 8'd10;
    sbox_10[164] = 8'd73;
    sbox_10[165] = 8'd6;
    sbox_10[166] = 8'd36;
    sbox_10[167] = 8'd92;
    sbox_10[168] = 8'd194;
    sbox_10[169] = 8'd211;
    sbox_10[170] = 8'd172;
    sbox_10[171] = 8'd98;
    sbox_10[172] = 8'd145;
    sbox_10[173] = 8'd149;
    sbox_10[174] = 8'd228;
    sbox_10[175] = 8'd121;
    sbox_10[176] = 8'd231;
    sbox_10[177] = 8'd200;
    sbox_10[178] = 8'd55;
    sbox_10[179] = 8'd109;
    sbox_10[180] = 8'd141;
    sbox_10[181] = 8'd213;
    sbox_10[182] = 8'd78;
    sbox_10[183] = 8'd169;
    sbox_10[184] = 8'd108;
    sbox_10[185] = 8'd86;
    sbox_10[186] = 8'd244;
    sbox_10[187] = 8'd234;
    sbox_10[188] = 8'd101;
    sbox_10[189] = 8'd122;
    sbox_10[190] = 8'd174;
    sbox_10[191] = 8'd8;
    sbox_10[192] = 8'd186;
    sbox_10[193] = 8'd120;
    sbox_10[194] = 8'd37;
    sbox_10[195] = 8'd46;
    sbox_10[196] = 8'd28;
    sbox_10[197] = 8'd166;
    sbox_10[198] = 8'd180;
    sbox_10[199] = 8'd198;
    sbox_10[200] = 8'd232;
    sbox_10[201] = 8'd221;
    sbox_10[202] = 8'd116;
    sbox_10[203] = 8'd31;
    sbox_10[204] = 8'd75;
    sbox_10[205] = 8'd189;
    sbox_10[206] = 8'd139;
    sbox_10[207] = 8'd138;
    sbox_10[208] = 8'd112;
    sbox_10[209] = 8'd62;
    sbox_10[210] = 8'd181;
    sbox_10[211] = 8'd102;
    sbox_10[212] = 8'd72;
    sbox_10[213] = 8'd3;
    sbox_10[214] = 8'd246;
    sbox_10[215] = 8'd14;
    sbox_10[216] = 8'd97;
    sbox_10[217] = 8'd53;
    sbox_10[218] = 8'd87;
    sbox_10[219] = 8'd185;
    sbox_10[220] = 8'd134;
    sbox_10[221] = 8'd193;
    sbox_10[222] = 8'd29;
    sbox_10[223] = 8'd158;
    sbox_10[224] = 8'd225;
    sbox_10[225] = 8'd248;
    sbox_10[226] = 8'd152;
    sbox_10[227] = 8'd17;
    sbox_10[228] = 8'd105;
    sbox_10[229] = 8'd217;
    sbox_10[230] = 8'd142;
    sbox_10[231] = 8'd148;
    sbox_10[232] = 8'd155;
    sbox_10[233] = 8'd30;
    sbox_10[234] = 8'd135;
    sbox_10[235] = 8'd233;
    sbox_10[236] = 8'd206;
    sbox_10[237] = 8'd85;
    sbox_10[238] = 8'd40;
    sbox_10[239] = 8'd223;
    sbox_10[240] = 8'd140;
    sbox_10[241] = 8'd161;
    sbox_10[242] = 8'd137;
    sbox_10[243] = 8'd13;
    sbox_10[244] = 8'd191;
    sbox_10[245] = 8'd230;
    sbox_10[246] = 8'd66;
    sbox_10[247] = 8'd104;
    sbox_10[248] = 8'd65;
    sbox_10[249] = 8'd153;
    sbox_10[250] = 8'd45;
    sbox_10[251] = 8'd15;
    sbox_10[252] = 8'd176;
    sbox_10[253] = 8'd84;
    sbox_10[254] = 8'd187;
    sbox_10[255] = 8'd22;
    sbox_11[0] = 8'd99;
    sbox_11[1] = 8'd124;
    sbox_11[2] = 8'd119;
    sbox_11[3] = 8'd123;
    sbox_11[4] = 8'd242;
    sbox_11[5] = 8'd107;
    sbox_11[6] = 8'd111;
    sbox_11[7] = 8'd197;
    sbox_11[8] = 8'd48;
    sbox_11[9] = 8'd1;
    sbox_11[10] = 8'd103;
    sbox_11[11] = 8'd43;
    sbox_11[12] = 8'd254;
    sbox_11[13] = 8'd215;
    sbox_11[14] = 8'd171;
    sbox_11[15] = 8'd118;
    sbox_11[16] = 8'd202;
    sbox_11[17] = 8'd130;
    sbox_11[18] = 8'd201;
    sbox_11[19] = 8'd125;
    sbox_11[20] = 8'd250;
    sbox_11[21] = 8'd89;
    sbox_11[22] = 8'd71;
    sbox_11[23] = 8'd240;
    sbox_11[24] = 8'd173;
    sbox_11[25] = 8'd212;
    sbox_11[26] = 8'd162;
    sbox_11[27] = 8'd175;
    sbox_11[28] = 8'd156;
    sbox_11[29] = 8'd164;
    sbox_11[30] = 8'd114;
    sbox_11[31] = 8'd192;
    sbox_11[32] = 8'd183;
    sbox_11[33] = 8'd253;
    sbox_11[34] = 8'd147;
    sbox_11[35] = 8'd38;
    sbox_11[36] = 8'd54;
    sbox_11[37] = 8'd63;
    sbox_11[38] = 8'd247;
    sbox_11[39] = 8'd204;
    sbox_11[40] = 8'd52;
    sbox_11[41] = 8'd165;
    sbox_11[42] = 8'd229;
    sbox_11[43] = 8'd241;
    sbox_11[44] = 8'd113;
    sbox_11[45] = 8'd216;
    sbox_11[46] = 8'd49;
    sbox_11[47] = 8'd21;
    sbox_11[48] = 8'd4;
    sbox_11[49] = 8'd199;
    sbox_11[50] = 8'd35;
    sbox_11[51] = 8'd195;
    sbox_11[52] = 8'd24;
    sbox_11[53] = 8'd150;
    sbox_11[54] = 8'd5;
    sbox_11[55] = 8'd154;
    sbox_11[56] = 8'd7;
    sbox_11[57] = 8'd18;
    sbox_11[58] = 8'd128;
    sbox_11[59] = 8'd226;
    sbox_11[60] = 8'd235;
    sbox_11[61] = 8'd39;
    sbox_11[62] = 8'd178;
    sbox_11[63] = 8'd117;
    sbox_11[64] = 8'd9;
    sbox_11[65] = 8'd131;
    sbox_11[66] = 8'd44;
    sbox_11[67] = 8'd26;
    sbox_11[68] = 8'd27;
    sbox_11[69] = 8'd110;
    sbox_11[70] = 8'd90;
    sbox_11[71] = 8'd160;
    sbox_11[72] = 8'd82;
    sbox_11[73] = 8'd59;
    sbox_11[74] = 8'd214;
    sbox_11[75] = 8'd179;
    sbox_11[76] = 8'd41;
    sbox_11[77] = 8'd227;
    sbox_11[78] = 8'd47;
    sbox_11[79] = 8'd132;
    sbox_11[80] = 8'd83;
    sbox_11[81] = 8'd209;
    sbox_11[82] = 8'd0;
    sbox_11[83] = 8'd237;
    sbox_11[84] = 8'd32;
    sbox_11[85] = 8'd252;
    sbox_11[86] = 8'd177;
    sbox_11[87] = 8'd91;
    sbox_11[88] = 8'd106;
    sbox_11[89] = 8'd203;
    sbox_11[90] = 8'd190;
    sbox_11[91] = 8'd57;
    sbox_11[92] = 8'd74;
    sbox_11[93] = 8'd76;
    sbox_11[94] = 8'd88;
    sbox_11[95] = 8'd207;
    sbox_11[96] = 8'd208;
    sbox_11[97] = 8'd239;
    sbox_11[98] = 8'd170;
    sbox_11[99] = 8'd251;
    sbox_11[100] = 8'd67;
    sbox_11[101] = 8'd77;
    sbox_11[102] = 8'd51;
    sbox_11[103] = 8'd133;
    sbox_11[104] = 8'd69;
    sbox_11[105] = 8'd249;
    sbox_11[106] = 8'd2;
    sbox_11[107] = 8'd127;
    sbox_11[108] = 8'd80;
    sbox_11[109] = 8'd60;
    sbox_11[110] = 8'd159;
    sbox_11[111] = 8'd168;
    sbox_11[112] = 8'd81;
    sbox_11[113] = 8'd163;
    sbox_11[114] = 8'd64;
    sbox_11[115] = 8'd143;
    sbox_11[116] = 8'd146;
    sbox_11[117] = 8'd157;
    sbox_11[118] = 8'd56;
    sbox_11[119] = 8'd245;
    sbox_11[120] = 8'd188;
    sbox_11[121] = 8'd182;
    sbox_11[122] = 8'd218;
    sbox_11[123] = 8'd33;
    sbox_11[124] = 8'd16;
    sbox_11[125] = 8'd255;
    sbox_11[126] = 8'd243;
    sbox_11[127] = 8'd210;
    sbox_11[128] = 8'd205;
    sbox_11[129] = 8'd12;
    sbox_11[130] = 8'd19;
    sbox_11[131] = 8'd236;
    sbox_11[132] = 8'd95;
    sbox_11[133] = 8'd151;
    sbox_11[134] = 8'd68;
    sbox_11[135] = 8'd23;
    sbox_11[136] = 8'd196;
    sbox_11[137] = 8'd167;
    sbox_11[138] = 8'd126;
    sbox_11[139] = 8'd61;
    sbox_11[140] = 8'd100;
    sbox_11[141] = 8'd93;
    sbox_11[142] = 8'd25;
    sbox_11[143] = 8'd115;
    sbox_11[144] = 8'd96;
    sbox_11[145] = 8'd129;
    sbox_11[146] = 8'd79;
    sbox_11[147] = 8'd220;
    sbox_11[148] = 8'd34;
    sbox_11[149] = 8'd42;
    sbox_11[150] = 8'd144;
    sbox_11[151] = 8'd136;
    sbox_11[152] = 8'd70;
    sbox_11[153] = 8'd238;
    sbox_11[154] = 8'd184;
    sbox_11[155] = 8'd20;
    sbox_11[156] = 8'd222;
    sbox_11[157] = 8'd94;
    sbox_11[158] = 8'd11;
    sbox_11[159] = 8'd219;
    sbox_11[160] = 8'd224;
    sbox_11[161] = 8'd50;
    sbox_11[162] = 8'd58;
    sbox_11[163] = 8'd10;
    sbox_11[164] = 8'd73;
    sbox_11[165] = 8'd6;
    sbox_11[166] = 8'd36;
    sbox_11[167] = 8'd92;
    sbox_11[168] = 8'd194;
    sbox_11[169] = 8'd211;
    sbox_11[170] = 8'd172;
    sbox_11[171] = 8'd98;
    sbox_11[172] = 8'd145;
    sbox_11[173] = 8'd149;
    sbox_11[174] = 8'd228;
    sbox_11[175] = 8'd121;
    sbox_11[176] = 8'd231;
    sbox_11[177] = 8'd200;
    sbox_11[178] = 8'd55;
    sbox_11[179] = 8'd109;
    sbox_11[180] = 8'd141;
    sbox_11[181] = 8'd213;
    sbox_11[182] = 8'd78;
    sbox_11[183] = 8'd169;
    sbox_11[184] = 8'd108;
    sbox_11[185] = 8'd86;
    sbox_11[186] = 8'd244;
    sbox_11[187] = 8'd234;
    sbox_11[188] = 8'd101;
    sbox_11[189] = 8'd122;
    sbox_11[190] = 8'd174;
    sbox_11[191] = 8'd8;
    sbox_11[192] = 8'd186;
    sbox_11[193] = 8'd120;
    sbox_11[194] = 8'd37;
    sbox_11[195] = 8'd46;
    sbox_11[196] = 8'd28;
    sbox_11[197] = 8'd166;
    sbox_11[198] = 8'd180;
    sbox_11[199] = 8'd198;
    sbox_11[200] = 8'd232;
    sbox_11[201] = 8'd221;
    sbox_11[202] = 8'd116;
    sbox_11[203] = 8'd31;
    sbox_11[204] = 8'd75;
    sbox_11[205] = 8'd189;
    sbox_11[206] = 8'd139;
    sbox_11[207] = 8'd138;
    sbox_11[208] = 8'd112;
    sbox_11[209] = 8'd62;
    sbox_11[210] = 8'd181;
    sbox_11[211] = 8'd102;
    sbox_11[212] = 8'd72;
    sbox_11[213] = 8'd3;
    sbox_11[214] = 8'd246;
    sbox_11[215] = 8'd14;
    sbox_11[216] = 8'd97;
    sbox_11[217] = 8'd53;
    sbox_11[218] = 8'd87;
    sbox_11[219] = 8'd185;
    sbox_11[220] = 8'd134;
    sbox_11[221] = 8'd193;
    sbox_11[222] = 8'd29;
    sbox_11[223] = 8'd158;
    sbox_11[224] = 8'd225;
    sbox_11[225] = 8'd248;
    sbox_11[226] = 8'd152;
    sbox_11[227] = 8'd17;
    sbox_11[228] = 8'd105;
    sbox_11[229] = 8'd217;
    sbox_11[230] = 8'd142;
    sbox_11[231] = 8'd148;
    sbox_11[232] = 8'd155;
    sbox_11[233] = 8'd30;
    sbox_11[234] = 8'd135;
    sbox_11[235] = 8'd233;
    sbox_11[236] = 8'd206;
    sbox_11[237] = 8'd85;
    sbox_11[238] = 8'd40;
    sbox_11[239] = 8'd223;
    sbox_11[240] = 8'd140;
    sbox_11[241] = 8'd161;
    sbox_11[242] = 8'd137;
    sbox_11[243] = 8'd13;
    sbox_11[244] = 8'd191;
    sbox_11[245] = 8'd230;
    sbox_11[246] = 8'd66;
    sbox_11[247] = 8'd104;
    sbox_11[248] = 8'd65;
    sbox_11[249] = 8'd153;
    sbox_11[250] = 8'd45;
    sbox_11[251] = 8'd15;
    sbox_11[252] = 8'd176;
    sbox_11[253] = 8'd84;
    sbox_11[254] = 8'd187;
    sbox_11[255] = 8'd22;
    sbox_12[0] = 8'd99;
    sbox_12[1] = 8'd124;
    sbox_12[2] = 8'd119;
    sbox_12[3] = 8'd123;
    sbox_12[4] = 8'd242;
    sbox_12[5] = 8'd107;
    sbox_12[6] = 8'd111;
    sbox_12[7] = 8'd197;
    sbox_12[8] = 8'd48;
    sbox_12[9] = 8'd1;
    sbox_12[10] = 8'd103;
    sbox_12[11] = 8'd43;
    sbox_12[12] = 8'd254;
    sbox_12[13] = 8'd215;
    sbox_12[14] = 8'd171;
    sbox_12[15] = 8'd118;
    sbox_12[16] = 8'd202;
    sbox_12[17] = 8'd130;
    sbox_12[18] = 8'd201;
    sbox_12[19] = 8'd125;
    sbox_12[20] = 8'd250;
    sbox_12[21] = 8'd89;
    sbox_12[22] = 8'd71;
    sbox_12[23] = 8'd240;
    sbox_12[24] = 8'd173;
    sbox_12[25] = 8'd212;
    sbox_12[26] = 8'd162;
    sbox_12[27] = 8'd175;
    sbox_12[28] = 8'd156;
    sbox_12[29] = 8'd164;
    sbox_12[30] = 8'd114;
    sbox_12[31] = 8'd192;
    sbox_12[32] = 8'd183;
    sbox_12[33] = 8'd253;
    sbox_12[34] = 8'd147;
    sbox_12[35] = 8'd38;
    sbox_12[36] = 8'd54;
    sbox_12[37] = 8'd63;
    sbox_12[38] = 8'd247;
    sbox_12[39] = 8'd204;
    sbox_12[40] = 8'd52;
    sbox_12[41] = 8'd165;
    sbox_12[42] = 8'd229;
    sbox_12[43] = 8'd241;
    sbox_12[44] = 8'd113;
    sbox_12[45] = 8'd216;
    sbox_12[46] = 8'd49;
    sbox_12[47] = 8'd21;
    sbox_12[48] = 8'd4;
    sbox_12[49] = 8'd199;
    sbox_12[50] = 8'd35;
    sbox_12[51] = 8'd195;
    sbox_12[52] = 8'd24;
    sbox_12[53] = 8'd150;
    sbox_12[54] = 8'd5;
    sbox_12[55] = 8'd154;
    sbox_12[56] = 8'd7;
    sbox_12[57] = 8'd18;
    sbox_12[58] = 8'd128;
    sbox_12[59] = 8'd226;
    sbox_12[60] = 8'd235;
    sbox_12[61] = 8'd39;
    sbox_12[62] = 8'd178;
    sbox_12[63] = 8'd117;
    sbox_12[64] = 8'd9;
    sbox_12[65] = 8'd131;
    sbox_12[66] = 8'd44;
    sbox_12[67] = 8'd26;
    sbox_12[68] = 8'd27;
    sbox_12[69] = 8'd110;
    sbox_12[70] = 8'd90;
    sbox_12[71] = 8'd160;
    sbox_12[72] = 8'd82;
    sbox_12[73] = 8'd59;
    sbox_12[74] = 8'd214;
    sbox_12[75] = 8'd179;
    sbox_12[76] = 8'd41;
    sbox_12[77] = 8'd227;
    sbox_12[78] = 8'd47;
    sbox_12[79] = 8'd132;
    sbox_12[80] = 8'd83;
    sbox_12[81] = 8'd209;
    sbox_12[82] = 8'd0;
    sbox_12[83] = 8'd237;
    sbox_12[84] = 8'd32;
    sbox_12[85] = 8'd252;
    sbox_12[86] = 8'd177;
    sbox_12[87] = 8'd91;
    sbox_12[88] = 8'd106;
    sbox_12[89] = 8'd203;
    sbox_12[90] = 8'd190;
    sbox_12[91] = 8'd57;
    sbox_12[92] = 8'd74;
    sbox_12[93] = 8'd76;
    sbox_12[94] = 8'd88;
    sbox_12[95] = 8'd207;
    sbox_12[96] = 8'd208;
    sbox_12[97] = 8'd239;
    sbox_12[98] = 8'd170;
    sbox_12[99] = 8'd251;
    sbox_12[100] = 8'd67;
    sbox_12[101] = 8'd77;
    sbox_12[102] = 8'd51;
    sbox_12[103] = 8'd133;
    sbox_12[104] = 8'd69;
    sbox_12[105] = 8'd249;
    sbox_12[106] = 8'd2;
    sbox_12[107] = 8'd127;
    sbox_12[108] = 8'd80;
    sbox_12[109] = 8'd60;
    sbox_12[110] = 8'd159;
    sbox_12[111] = 8'd168;
    sbox_12[112] = 8'd81;
    sbox_12[113] = 8'd163;
    sbox_12[114] = 8'd64;
    sbox_12[115] = 8'd143;
    sbox_12[116] = 8'd146;
    sbox_12[117] = 8'd157;
    sbox_12[118] = 8'd56;
    sbox_12[119] = 8'd245;
    sbox_12[120] = 8'd188;
    sbox_12[121] = 8'd182;
    sbox_12[122] = 8'd218;
    sbox_12[123] = 8'd33;
    sbox_12[124] = 8'd16;
    sbox_12[125] = 8'd255;
    sbox_12[126] = 8'd243;
    sbox_12[127] = 8'd210;
    sbox_12[128] = 8'd205;
    sbox_12[129] = 8'd12;
    sbox_12[130] = 8'd19;
    sbox_12[131] = 8'd236;
    sbox_12[132] = 8'd95;
    sbox_12[133] = 8'd151;
    sbox_12[134] = 8'd68;
    sbox_12[135] = 8'd23;
    sbox_12[136] = 8'd196;
    sbox_12[137] = 8'd167;
    sbox_12[138] = 8'd126;
    sbox_12[139] = 8'd61;
    sbox_12[140] = 8'd100;
    sbox_12[141] = 8'd93;
    sbox_12[142] = 8'd25;
    sbox_12[143] = 8'd115;
    sbox_12[144] = 8'd96;
    sbox_12[145] = 8'd129;
    sbox_12[146] = 8'd79;
    sbox_12[147] = 8'd220;
    sbox_12[148] = 8'd34;
    sbox_12[149] = 8'd42;
    sbox_12[150] = 8'd144;
    sbox_12[151] = 8'd136;
    sbox_12[152] = 8'd70;
    sbox_12[153] = 8'd238;
    sbox_12[154] = 8'd184;
    sbox_12[155] = 8'd20;
    sbox_12[156] = 8'd222;
    sbox_12[157] = 8'd94;
    sbox_12[158] = 8'd11;
    sbox_12[159] = 8'd219;
    sbox_12[160] = 8'd224;
    sbox_12[161] = 8'd50;
    sbox_12[162] = 8'd58;
    sbox_12[163] = 8'd10;
    sbox_12[164] = 8'd73;
    sbox_12[165] = 8'd6;
    sbox_12[166] = 8'd36;
    sbox_12[167] = 8'd92;
    sbox_12[168] = 8'd194;
    sbox_12[169] = 8'd211;
    sbox_12[170] = 8'd172;
    sbox_12[171] = 8'd98;
    sbox_12[172] = 8'd145;
    sbox_12[173] = 8'd149;
    sbox_12[174] = 8'd228;
    sbox_12[175] = 8'd121;
    sbox_12[176] = 8'd231;
    sbox_12[177] = 8'd200;
    sbox_12[178] = 8'd55;
    sbox_12[179] = 8'd109;
    sbox_12[180] = 8'd141;
    sbox_12[181] = 8'd213;
    sbox_12[182] = 8'd78;
    sbox_12[183] = 8'd169;
    sbox_12[184] = 8'd108;
    sbox_12[185] = 8'd86;
    sbox_12[186] = 8'd244;
    sbox_12[187] = 8'd234;
    sbox_12[188] = 8'd101;
    sbox_12[189] = 8'd122;
    sbox_12[190] = 8'd174;
    sbox_12[191] = 8'd8;
    sbox_12[192] = 8'd186;
    sbox_12[193] = 8'd120;
    sbox_12[194] = 8'd37;
    sbox_12[195] = 8'd46;
    sbox_12[196] = 8'd28;
    sbox_12[197] = 8'd166;
    sbox_12[198] = 8'd180;
    sbox_12[199] = 8'd198;
    sbox_12[200] = 8'd232;
    sbox_12[201] = 8'd221;
    sbox_12[202] = 8'd116;
    sbox_12[203] = 8'd31;
    sbox_12[204] = 8'd75;
    sbox_12[205] = 8'd189;
    sbox_12[206] = 8'd139;
    sbox_12[207] = 8'd138;
    sbox_12[208] = 8'd112;
    sbox_12[209] = 8'd62;
    sbox_12[210] = 8'd181;
    sbox_12[211] = 8'd102;
    sbox_12[212] = 8'd72;
    sbox_12[213] = 8'd3;
    sbox_12[214] = 8'd246;
    sbox_12[215] = 8'd14;
    sbox_12[216] = 8'd97;
    sbox_12[217] = 8'd53;
    sbox_12[218] = 8'd87;
    sbox_12[219] = 8'd185;
    sbox_12[220] = 8'd134;
    sbox_12[221] = 8'd193;
    sbox_12[222] = 8'd29;
    sbox_12[223] = 8'd158;
    sbox_12[224] = 8'd225;
    sbox_12[225] = 8'd248;
    sbox_12[226] = 8'd152;
    sbox_12[227] = 8'd17;
    sbox_12[228] = 8'd105;
    sbox_12[229] = 8'd217;
    sbox_12[230] = 8'd142;
    sbox_12[231] = 8'd148;
    sbox_12[232] = 8'd155;
    sbox_12[233] = 8'd30;
    sbox_12[234] = 8'd135;
    sbox_12[235] = 8'd233;
    sbox_12[236] = 8'd206;
    sbox_12[237] = 8'd85;
    sbox_12[238] = 8'd40;
    sbox_12[239] = 8'd223;
    sbox_12[240] = 8'd140;
    sbox_12[241] = 8'd161;
    sbox_12[242] = 8'd137;
    sbox_12[243] = 8'd13;
    sbox_12[244] = 8'd191;
    sbox_12[245] = 8'd230;
    sbox_12[246] = 8'd66;
    sbox_12[247] = 8'd104;
    sbox_12[248] = 8'd65;
    sbox_12[249] = 8'd153;
    sbox_12[250] = 8'd45;
    sbox_12[251] = 8'd15;
    sbox_12[252] = 8'd176;
    sbox_12[253] = 8'd84;
    sbox_12[254] = 8'd187;
    sbox_12[255] = 8'd22;
    sbox_13[0] = 8'd99;
    sbox_13[1] = 8'd124;
    sbox_13[2] = 8'd119;
    sbox_13[3] = 8'd123;
    sbox_13[4] = 8'd242;
    sbox_13[5] = 8'd107;
    sbox_13[6] = 8'd111;
    sbox_13[7] = 8'd197;
    sbox_13[8] = 8'd48;
    sbox_13[9] = 8'd1;
    sbox_13[10] = 8'd103;
    sbox_13[11] = 8'd43;
    sbox_13[12] = 8'd254;
    sbox_13[13] = 8'd215;
    sbox_13[14] = 8'd171;
    sbox_13[15] = 8'd118;
    sbox_13[16] = 8'd202;
    sbox_13[17] = 8'd130;
    sbox_13[18] = 8'd201;
    sbox_13[19] = 8'd125;
    sbox_13[20] = 8'd250;
    sbox_13[21] = 8'd89;
    sbox_13[22] = 8'd71;
    sbox_13[23] = 8'd240;
    sbox_13[24] = 8'd173;
    sbox_13[25] = 8'd212;
    sbox_13[26] = 8'd162;
    sbox_13[27] = 8'd175;
    sbox_13[28] = 8'd156;
    sbox_13[29] = 8'd164;
    sbox_13[30] = 8'd114;
    sbox_13[31] = 8'd192;
    sbox_13[32] = 8'd183;
    sbox_13[33] = 8'd253;
    sbox_13[34] = 8'd147;
    sbox_13[35] = 8'd38;
    sbox_13[36] = 8'd54;
    sbox_13[37] = 8'd63;
    sbox_13[38] = 8'd247;
    sbox_13[39] = 8'd204;
    sbox_13[40] = 8'd52;
    sbox_13[41] = 8'd165;
    sbox_13[42] = 8'd229;
    sbox_13[43] = 8'd241;
    sbox_13[44] = 8'd113;
    sbox_13[45] = 8'd216;
    sbox_13[46] = 8'd49;
    sbox_13[47] = 8'd21;
    sbox_13[48] = 8'd4;
    sbox_13[49] = 8'd199;
    sbox_13[50] = 8'd35;
    sbox_13[51] = 8'd195;
    sbox_13[52] = 8'd24;
    sbox_13[53] = 8'd150;
    sbox_13[54] = 8'd5;
    sbox_13[55] = 8'd154;
    sbox_13[56] = 8'd7;
    sbox_13[57] = 8'd18;
    sbox_13[58] = 8'd128;
    sbox_13[59] = 8'd226;
    sbox_13[60] = 8'd235;
    sbox_13[61] = 8'd39;
    sbox_13[62] = 8'd178;
    sbox_13[63] = 8'd117;
    sbox_13[64] = 8'd9;
    sbox_13[65] = 8'd131;
    sbox_13[66] = 8'd44;
    sbox_13[67] = 8'd26;
    sbox_13[68] = 8'd27;
    sbox_13[69] = 8'd110;
    sbox_13[70] = 8'd90;
    sbox_13[71] = 8'd160;
    sbox_13[72] = 8'd82;
    sbox_13[73] = 8'd59;
    sbox_13[74] = 8'd214;
    sbox_13[75] = 8'd179;
    sbox_13[76] = 8'd41;
    sbox_13[77] = 8'd227;
    sbox_13[78] = 8'd47;
    sbox_13[79] = 8'd132;
    sbox_13[80] = 8'd83;
    sbox_13[81] = 8'd209;
    sbox_13[82] = 8'd0;
    sbox_13[83] = 8'd237;
    sbox_13[84] = 8'd32;
    sbox_13[85] = 8'd252;
    sbox_13[86] = 8'd177;
    sbox_13[87] = 8'd91;
    sbox_13[88] = 8'd106;
    sbox_13[89] = 8'd203;
    sbox_13[90] = 8'd190;
    sbox_13[91] = 8'd57;
    sbox_13[92] = 8'd74;
    sbox_13[93] = 8'd76;
    sbox_13[94] = 8'd88;
    sbox_13[95] = 8'd207;
    sbox_13[96] = 8'd208;
    sbox_13[97] = 8'd239;
    sbox_13[98] = 8'd170;
    sbox_13[99] = 8'd251;
    sbox_13[100] = 8'd67;
    sbox_13[101] = 8'd77;
    sbox_13[102] = 8'd51;
    sbox_13[103] = 8'd133;
    sbox_13[104] = 8'd69;
    sbox_13[105] = 8'd249;
    sbox_13[106] = 8'd2;
    sbox_13[107] = 8'd127;
    sbox_13[108] = 8'd80;
    sbox_13[109] = 8'd60;
    sbox_13[110] = 8'd159;
    sbox_13[111] = 8'd168;
    sbox_13[112] = 8'd81;
    sbox_13[113] = 8'd163;
    sbox_13[114] = 8'd64;
    sbox_13[115] = 8'd143;
    sbox_13[116] = 8'd146;
    sbox_13[117] = 8'd157;
    sbox_13[118] = 8'd56;
    sbox_13[119] = 8'd245;
    sbox_13[120] = 8'd188;
    sbox_13[121] = 8'd182;
    sbox_13[122] = 8'd218;
    sbox_13[123] = 8'd33;
    sbox_13[124] = 8'd16;
    sbox_13[125] = 8'd255;
    sbox_13[126] = 8'd243;
    sbox_13[127] = 8'd210;
    sbox_13[128] = 8'd205;
    sbox_13[129] = 8'd12;
    sbox_13[130] = 8'd19;
    sbox_13[131] = 8'd236;
    sbox_13[132] = 8'd95;
    sbox_13[133] = 8'd151;
    sbox_13[134] = 8'd68;
    sbox_13[135] = 8'd23;
    sbox_13[136] = 8'd196;
    sbox_13[137] = 8'd167;
    sbox_13[138] = 8'd126;
    sbox_13[139] = 8'd61;
    sbox_13[140] = 8'd100;
    sbox_13[141] = 8'd93;
    sbox_13[142] = 8'd25;
    sbox_13[143] = 8'd115;
    sbox_13[144] = 8'd96;
    sbox_13[145] = 8'd129;
    sbox_13[146] = 8'd79;
    sbox_13[147] = 8'd220;
    sbox_13[148] = 8'd34;
    sbox_13[149] = 8'd42;
    sbox_13[150] = 8'd144;
    sbox_13[151] = 8'd136;
    sbox_13[152] = 8'd70;
    sbox_13[153] = 8'd238;
    sbox_13[154] = 8'd184;
    sbox_13[155] = 8'd20;
    sbox_13[156] = 8'd222;
    sbox_13[157] = 8'd94;
    sbox_13[158] = 8'd11;
    sbox_13[159] = 8'd219;
    sbox_13[160] = 8'd224;
    sbox_13[161] = 8'd50;
    sbox_13[162] = 8'd58;
    sbox_13[163] = 8'd10;
    sbox_13[164] = 8'd73;
    sbox_13[165] = 8'd6;
    sbox_13[166] = 8'd36;
    sbox_13[167] = 8'd92;
    sbox_13[168] = 8'd194;
    sbox_13[169] = 8'd211;
    sbox_13[170] = 8'd172;
    sbox_13[171] = 8'd98;
    sbox_13[172] = 8'd145;
    sbox_13[173] = 8'd149;
    sbox_13[174] = 8'd228;
    sbox_13[175] = 8'd121;
    sbox_13[176] = 8'd231;
    sbox_13[177] = 8'd200;
    sbox_13[178] = 8'd55;
    sbox_13[179] = 8'd109;
    sbox_13[180] = 8'd141;
    sbox_13[181] = 8'd213;
    sbox_13[182] = 8'd78;
    sbox_13[183] = 8'd169;
    sbox_13[184] = 8'd108;
    sbox_13[185] = 8'd86;
    sbox_13[186] = 8'd244;
    sbox_13[187] = 8'd234;
    sbox_13[188] = 8'd101;
    sbox_13[189] = 8'd122;
    sbox_13[190] = 8'd174;
    sbox_13[191] = 8'd8;
    sbox_13[192] = 8'd186;
    sbox_13[193] = 8'd120;
    sbox_13[194] = 8'd37;
    sbox_13[195] = 8'd46;
    sbox_13[196] = 8'd28;
    sbox_13[197] = 8'd166;
    sbox_13[198] = 8'd180;
    sbox_13[199] = 8'd198;
    sbox_13[200] = 8'd232;
    sbox_13[201] = 8'd221;
    sbox_13[202] = 8'd116;
    sbox_13[203] = 8'd31;
    sbox_13[204] = 8'd75;
    sbox_13[205] = 8'd189;
    sbox_13[206] = 8'd139;
    sbox_13[207] = 8'd138;
    sbox_13[208] = 8'd112;
    sbox_13[209] = 8'd62;
    sbox_13[210] = 8'd181;
    sbox_13[211] = 8'd102;
    sbox_13[212] = 8'd72;
    sbox_13[213] = 8'd3;
    sbox_13[214] = 8'd246;
    sbox_13[215] = 8'd14;
    sbox_13[216] = 8'd97;
    sbox_13[217] = 8'd53;
    sbox_13[218] = 8'd87;
    sbox_13[219] = 8'd185;
    sbox_13[220] = 8'd134;
    sbox_13[221] = 8'd193;
    sbox_13[222] = 8'd29;
    sbox_13[223] = 8'd158;
    sbox_13[224] = 8'd225;
    sbox_13[225] = 8'd248;
    sbox_13[226] = 8'd152;
    sbox_13[227] = 8'd17;
    sbox_13[228] = 8'd105;
    sbox_13[229] = 8'd217;
    sbox_13[230] = 8'd142;
    sbox_13[231] = 8'd148;
    sbox_13[232] = 8'd155;
    sbox_13[233] = 8'd30;
    sbox_13[234] = 8'd135;
    sbox_13[235] = 8'd233;
    sbox_13[236] = 8'd206;
    sbox_13[237] = 8'd85;
    sbox_13[238] = 8'd40;
    sbox_13[239] = 8'd223;
    sbox_13[240] = 8'd140;
    sbox_13[241] = 8'd161;
    sbox_13[242] = 8'd137;
    sbox_13[243] = 8'd13;
    sbox_13[244] = 8'd191;
    sbox_13[245] = 8'd230;
    sbox_13[246] = 8'd66;
    sbox_13[247] = 8'd104;
    sbox_13[248] = 8'd65;
    sbox_13[249] = 8'd153;
    sbox_13[250] = 8'd45;
    sbox_13[251] = 8'd15;
    sbox_13[252] = 8'd176;
    sbox_13[253] = 8'd84;
    sbox_13[254] = 8'd187;
    sbox_13[255] = 8'd22;
    sbox_14[0] = 8'd99;
    sbox_14[1] = 8'd124;
    sbox_14[2] = 8'd119;
    sbox_14[3] = 8'd123;
    sbox_14[4] = 8'd242;
    sbox_14[5] = 8'd107;
    sbox_14[6] = 8'd111;
    sbox_14[7] = 8'd197;
    sbox_14[8] = 8'd48;
    sbox_14[9] = 8'd1;
    sbox_14[10] = 8'd103;
    sbox_14[11] = 8'd43;
    sbox_14[12] = 8'd254;
    sbox_14[13] = 8'd215;
    sbox_14[14] = 8'd171;
    sbox_14[15] = 8'd118;
    sbox_14[16] = 8'd202;
    sbox_14[17] = 8'd130;
    sbox_14[18] = 8'd201;
    sbox_14[19] = 8'd125;
    sbox_14[20] = 8'd250;
    sbox_14[21] = 8'd89;
    sbox_14[22] = 8'd71;
    sbox_14[23] = 8'd240;
    sbox_14[24] = 8'd173;
    sbox_14[25] = 8'd212;
    sbox_14[26] = 8'd162;
    sbox_14[27] = 8'd175;
    sbox_14[28] = 8'd156;
    sbox_14[29] = 8'd164;
    sbox_14[30] = 8'd114;
    sbox_14[31] = 8'd192;
    sbox_14[32] = 8'd183;
    sbox_14[33] = 8'd253;
    sbox_14[34] = 8'd147;
    sbox_14[35] = 8'd38;
    sbox_14[36] = 8'd54;
    sbox_14[37] = 8'd63;
    sbox_14[38] = 8'd247;
    sbox_14[39] = 8'd204;
    sbox_14[40] = 8'd52;
    sbox_14[41] = 8'd165;
    sbox_14[42] = 8'd229;
    sbox_14[43] = 8'd241;
    sbox_14[44] = 8'd113;
    sbox_14[45] = 8'd216;
    sbox_14[46] = 8'd49;
    sbox_14[47] = 8'd21;
    sbox_14[48] = 8'd4;
    sbox_14[49] = 8'd199;
    sbox_14[50] = 8'd35;
    sbox_14[51] = 8'd195;
    sbox_14[52] = 8'd24;
    sbox_14[53] = 8'd150;
    sbox_14[54] = 8'd5;
    sbox_14[55] = 8'd154;
    sbox_14[56] = 8'd7;
    sbox_14[57] = 8'd18;
    sbox_14[58] = 8'd128;
    sbox_14[59] = 8'd226;
    sbox_14[60] = 8'd235;
    sbox_14[61] = 8'd39;
    sbox_14[62] = 8'd178;
    sbox_14[63] = 8'd117;
    sbox_14[64] = 8'd9;
    sbox_14[65] = 8'd131;
    sbox_14[66] = 8'd44;
    sbox_14[67] = 8'd26;
    sbox_14[68] = 8'd27;
    sbox_14[69] = 8'd110;
    sbox_14[70] = 8'd90;
    sbox_14[71] = 8'd160;
    sbox_14[72] = 8'd82;
    sbox_14[73] = 8'd59;
    sbox_14[74] = 8'd214;
    sbox_14[75] = 8'd179;
    sbox_14[76] = 8'd41;
    sbox_14[77] = 8'd227;
    sbox_14[78] = 8'd47;
    sbox_14[79] = 8'd132;
    sbox_14[80] = 8'd83;
    sbox_14[81] = 8'd209;
    sbox_14[82] = 8'd0;
    sbox_14[83] = 8'd237;
    sbox_14[84] = 8'd32;
    sbox_14[85] = 8'd252;
    sbox_14[86] = 8'd177;
    sbox_14[87] = 8'd91;
    sbox_14[88] = 8'd106;
    sbox_14[89] = 8'd203;
    sbox_14[90] = 8'd190;
    sbox_14[91] = 8'd57;
    sbox_14[92] = 8'd74;
    sbox_14[93] = 8'd76;
    sbox_14[94] = 8'd88;
    sbox_14[95] = 8'd207;
    sbox_14[96] = 8'd208;
    sbox_14[97] = 8'd239;
    sbox_14[98] = 8'd170;
    sbox_14[99] = 8'd251;
    sbox_14[100] = 8'd67;
    sbox_14[101] = 8'd77;
    sbox_14[102] = 8'd51;
    sbox_14[103] = 8'd133;
    sbox_14[104] = 8'd69;
    sbox_14[105] = 8'd249;
    sbox_14[106] = 8'd2;
    sbox_14[107] = 8'd127;
    sbox_14[108] = 8'd80;
    sbox_14[109] = 8'd60;
    sbox_14[110] = 8'd159;
    sbox_14[111] = 8'd168;
    sbox_14[112] = 8'd81;
    sbox_14[113] = 8'd163;
    sbox_14[114] = 8'd64;
    sbox_14[115] = 8'd143;
    sbox_14[116] = 8'd146;
    sbox_14[117] = 8'd157;
    sbox_14[118] = 8'd56;
    sbox_14[119] = 8'd245;
    sbox_14[120] = 8'd188;
    sbox_14[121] = 8'd182;
    sbox_14[122] = 8'd218;
    sbox_14[123] = 8'd33;
    sbox_14[124] = 8'd16;
    sbox_14[125] = 8'd255;
    sbox_14[126] = 8'd243;
    sbox_14[127] = 8'd210;
    sbox_14[128] = 8'd205;
    sbox_14[129] = 8'd12;
    sbox_14[130] = 8'd19;
    sbox_14[131] = 8'd236;
    sbox_14[132] = 8'd95;
    sbox_14[133] = 8'd151;
    sbox_14[134] = 8'd68;
    sbox_14[135] = 8'd23;
    sbox_14[136] = 8'd196;
    sbox_14[137] = 8'd167;
    sbox_14[138] = 8'd126;
    sbox_14[139] = 8'd61;
    sbox_14[140] = 8'd100;
    sbox_14[141] = 8'd93;
    sbox_14[142] = 8'd25;
    sbox_14[143] = 8'd115;
    sbox_14[144] = 8'd96;
    sbox_14[145] = 8'd129;
    sbox_14[146] = 8'd79;
    sbox_14[147] = 8'd220;
    sbox_14[148] = 8'd34;
    sbox_14[149] = 8'd42;
    sbox_14[150] = 8'd144;
    sbox_14[151] = 8'd136;
    sbox_14[152] = 8'd70;
    sbox_14[153] = 8'd238;
    sbox_14[154] = 8'd184;
    sbox_14[155] = 8'd20;
    sbox_14[156] = 8'd222;
    sbox_14[157] = 8'd94;
    sbox_14[158] = 8'd11;
    sbox_14[159] = 8'd219;
    sbox_14[160] = 8'd224;
    sbox_14[161] = 8'd50;
    sbox_14[162] = 8'd58;
    sbox_14[163] = 8'd10;
    sbox_14[164] = 8'd73;
    sbox_14[165] = 8'd6;
    sbox_14[166] = 8'd36;
    sbox_14[167] = 8'd92;
    sbox_14[168] = 8'd194;
    sbox_14[169] = 8'd211;
    sbox_14[170] = 8'd172;
    sbox_14[171] = 8'd98;
    sbox_14[172] = 8'd145;
    sbox_14[173] = 8'd149;
    sbox_14[174] = 8'd228;
    sbox_14[175] = 8'd121;
    sbox_14[176] = 8'd231;
    sbox_14[177] = 8'd200;
    sbox_14[178] = 8'd55;
    sbox_14[179] = 8'd109;
    sbox_14[180] = 8'd141;
    sbox_14[181] = 8'd213;
    sbox_14[182] = 8'd78;
    sbox_14[183] = 8'd169;
    sbox_14[184] = 8'd108;
    sbox_14[185] = 8'd86;
    sbox_14[186] = 8'd244;
    sbox_14[187] = 8'd234;
    sbox_14[188] = 8'd101;
    sbox_14[189] = 8'd122;
    sbox_14[190] = 8'd174;
    sbox_14[191] = 8'd8;
    sbox_14[192] = 8'd186;
    sbox_14[193] = 8'd120;
    sbox_14[194] = 8'd37;
    sbox_14[195] = 8'd46;
    sbox_14[196] = 8'd28;
    sbox_14[197] = 8'd166;
    sbox_14[198] = 8'd180;
    sbox_14[199] = 8'd198;
    sbox_14[200] = 8'd232;
    sbox_14[201] = 8'd221;
    sbox_14[202] = 8'd116;
    sbox_14[203] = 8'd31;
    sbox_14[204] = 8'd75;
    sbox_14[205] = 8'd189;
    sbox_14[206] = 8'd139;
    sbox_14[207] = 8'd138;
    sbox_14[208] = 8'd112;
    sbox_14[209] = 8'd62;
    sbox_14[210] = 8'd181;
    sbox_14[211] = 8'd102;
    sbox_14[212] = 8'd72;
    sbox_14[213] = 8'd3;
    sbox_14[214] = 8'd246;
    sbox_14[215] = 8'd14;
    sbox_14[216] = 8'd97;
    sbox_14[217] = 8'd53;
    sbox_14[218] = 8'd87;
    sbox_14[219] = 8'd185;
    sbox_14[220] = 8'd134;
    sbox_14[221] = 8'd193;
    sbox_14[222] = 8'd29;
    sbox_14[223] = 8'd158;
    sbox_14[224] = 8'd225;
    sbox_14[225] = 8'd248;
    sbox_14[226] = 8'd152;
    sbox_14[227] = 8'd17;
    sbox_14[228] = 8'd105;
    sbox_14[229] = 8'd217;
    sbox_14[230] = 8'd142;
    sbox_14[231] = 8'd148;
    sbox_14[232] = 8'd155;
    sbox_14[233] = 8'd30;
    sbox_14[234] = 8'd135;
    sbox_14[235] = 8'd233;
    sbox_14[236] = 8'd206;
    sbox_14[237] = 8'd85;
    sbox_14[238] = 8'd40;
    sbox_14[239] = 8'd223;
    sbox_14[240] = 8'd140;
    sbox_14[241] = 8'd161;
    sbox_14[242] = 8'd137;
    sbox_14[243] = 8'd13;
    sbox_14[244] = 8'd191;
    sbox_14[245] = 8'd230;
    sbox_14[246] = 8'd66;
    sbox_14[247] = 8'd104;
    sbox_14[248] = 8'd65;
    sbox_14[249] = 8'd153;
    sbox_14[250] = 8'd45;
    sbox_14[251] = 8'd15;
    sbox_14[252] = 8'd176;
    sbox_14[253] = 8'd84;
    sbox_14[254] = 8'd187;
    sbox_14[255] = 8'd22;
    sbox_15[0] = 8'd99;
    sbox_15[1] = 8'd124;
    sbox_15[2] = 8'd119;
    sbox_15[3] = 8'd123;
    sbox_15[4] = 8'd242;
    sbox_15[5] = 8'd107;
    sbox_15[6] = 8'd111;
    sbox_15[7] = 8'd197;
    sbox_15[8] = 8'd48;
    sbox_15[9] = 8'd1;
    sbox_15[10] = 8'd103;
    sbox_15[11] = 8'd43;
    sbox_15[12] = 8'd254;
    sbox_15[13] = 8'd215;
    sbox_15[14] = 8'd171;
    sbox_15[15] = 8'd118;
    sbox_15[16] = 8'd202;
    sbox_15[17] = 8'd130;
    sbox_15[18] = 8'd201;
    sbox_15[19] = 8'd125;
    sbox_15[20] = 8'd250;
    sbox_15[21] = 8'd89;
    sbox_15[22] = 8'd71;
    sbox_15[23] = 8'd240;
    sbox_15[24] = 8'd173;
    sbox_15[25] = 8'd212;
    sbox_15[26] = 8'd162;
    sbox_15[27] = 8'd175;
    sbox_15[28] = 8'd156;
    sbox_15[29] = 8'd164;
    sbox_15[30] = 8'd114;
    sbox_15[31] = 8'd192;
    sbox_15[32] = 8'd183;
    sbox_15[33] = 8'd253;
    sbox_15[34] = 8'd147;
    sbox_15[35] = 8'd38;
    sbox_15[36] = 8'd54;
    sbox_15[37] = 8'd63;
    sbox_15[38] = 8'd247;
    sbox_15[39] = 8'd204;
    sbox_15[40] = 8'd52;
    sbox_15[41] = 8'd165;
    sbox_15[42] = 8'd229;
    sbox_15[43] = 8'd241;
    sbox_15[44] = 8'd113;
    sbox_15[45] = 8'd216;
    sbox_15[46] = 8'd49;
    sbox_15[47] = 8'd21;
    sbox_15[48] = 8'd4;
    sbox_15[49] = 8'd199;
    sbox_15[50] = 8'd35;
    sbox_15[51] = 8'd195;
    sbox_15[52] = 8'd24;
    sbox_15[53] = 8'd150;
    sbox_15[54] = 8'd5;
    sbox_15[55] = 8'd154;
    sbox_15[56] = 8'd7;
    sbox_15[57] = 8'd18;
    sbox_15[58] = 8'd128;
    sbox_15[59] = 8'd226;
    sbox_15[60] = 8'd235;
    sbox_15[61] = 8'd39;
    sbox_15[62] = 8'd178;
    sbox_15[63] = 8'd117;
    sbox_15[64] = 8'd9;
    sbox_15[65] = 8'd131;
    sbox_15[66] = 8'd44;
    sbox_15[67] = 8'd26;
    sbox_15[68] = 8'd27;
    sbox_15[69] = 8'd110;
    sbox_15[70] = 8'd90;
    sbox_15[71] = 8'd160;
    sbox_15[72] = 8'd82;
    sbox_15[73] = 8'd59;
    sbox_15[74] = 8'd214;
    sbox_15[75] = 8'd179;
    sbox_15[76] = 8'd41;
    sbox_15[77] = 8'd227;
    sbox_15[78] = 8'd47;
    sbox_15[79] = 8'd132;
    sbox_15[80] = 8'd83;
    sbox_15[81] = 8'd209;
    sbox_15[82] = 8'd0;
    sbox_15[83] = 8'd237;
    sbox_15[84] = 8'd32;
    sbox_15[85] = 8'd252;
    sbox_15[86] = 8'd177;
    sbox_15[87] = 8'd91;
    sbox_15[88] = 8'd106;
    sbox_15[89] = 8'd203;
    sbox_15[90] = 8'd190;
    sbox_15[91] = 8'd57;
    sbox_15[92] = 8'd74;
    sbox_15[93] = 8'd76;
    sbox_15[94] = 8'd88;
    sbox_15[95] = 8'd207;
    sbox_15[96] = 8'd208;
    sbox_15[97] = 8'd239;
    sbox_15[98] = 8'd170;
    sbox_15[99] = 8'd251;
    sbox_15[100] = 8'd67;
    sbox_15[101] = 8'd77;
    sbox_15[102] = 8'd51;
    sbox_15[103] = 8'd133;
    sbox_15[104] = 8'd69;
    sbox_15[105] = 8'd249;
    sbox_15[106] = 8'd2;
    sbox_15[107] = 8'd127;
    sbox_15[108] = 8'd80;
    sbox_15[109] = 8'd60;
    sbox_15[110] = 8'd159;
    sbox_15[111] = 8'd168;
    sbox_15[112] = 8'd81;
    sbox_15[113] = 8'd163;
    sbox_15[114] = 8'd64;
    sbox_15[115] = 8'd143;
    sbox_15[116] = 8'd146;
    sbox_15[117] = 8'd157;
    sbox_15[118] = 8'd56;
    sbox_15[119] = 8'd245;
    sbox_15[120] = 8'd188;
    sbox_15[121] = 8'd182;
    sbox_15[122] = 8'd218;
    sbox_15[123] = 8'd33;
    sbox_15[124] = 8'd16;
    sbox_15[125] = 8'd255;
    sbox_15[126] = 8'd243;
    sbox_15[127] = 8'd210;
    sbox_15[128] = 8'd205;
    sbox_15[129] = 8'd12;
    sbox_15[130] = 8'd19;
    sbox_15[131] = 8'd236;
    sbox_15[132] = 8'd95;
    sbox_15[133] = 8'd151;
    sbox_15[134] = 8'd68;
    sbox_15[135] = 8'd23;
    sbox_15[136] = 8'd196;
    sbox_15[137] = 8'd167;
    sbox_15[138] = 8'd126;
    sbox_15[139] = 8'd61;
    sbox_15[140] = 8'd100;
    sbox_15[141] = 8'd93;
    sbox_15[142] = 8'd25;
    sbox_15[143] = 8'd115;
    sbox_15[144] = 8'd96;
    sbox_15[145] = 8'd129;
    sbox_15[146] = 8'd79;
    sbox_15[147] = 8'd220;
    sbox_15[148] = 8'd34;
    sbox_15[149] = 8'd42;
    sbox_15[150] = 8'd144;
    sbox_15[151] = 8'd136;
    sbox_15[152] = 8'd70;
    sbox_15[153] = 8'd238;
    sbox_15[154] = 8'd184;
    sbox_15[155] = 8'd20;
    sbox_15[156] = 8'd222;
    sbox_15[157] = 8'd94;
    sbox_15[158] = 8'd11;
    sbox_15[159] = 8'd219;
    sbox_15[160] = 8'd224;
    sbox_15[161] = 8'd50;
    sbox_15[162] = 8'd58;
    sbox_15[163] = 8'd10;
    sbox_15[164] = 8'd73;
    sbox_15[165] = 8'd6;
    sbox_15[166] = 8'd36;
    sbox_15[167] = 8'd92;
    sbox_15[168] = 8'd194;
    sbox_15[169] = 8'd211;
    sbox_15[170] = 8'd172;
    sbox_15[171] = 8'd98;
    sbox_15[172] = 8'd145;
    sbox_15[173] = 8'd149;
    sbox_15[174] = 8'd228;
    sbox_15[175] = 8'd121;
    sbox_15[176] = 8'd231;
    sbox_15[177] = 8'd200;
    sbox_15[178] = 8'd55;
    sbox_15[179] = 8'd109;
    sbox_15[180] = 8'd141;
    sbox_15[181] = 8'd213;
    sbox_15[182] = 8'd78;
    sbox_15[183] = 8'd169;
    sbox_15[184] = 8'd108;
    sbox_15[185] = 8'd86;
    sbox_15[186] = 8'd244;
    sbox_15[187] = 8'd234;
    sbox_15[188] = 8'd101;
    sbox_15[189] = 8'd122;
    sbox_15[190] = 8'd174;
    sbox_15[191] = 8'd8;
    sbox_15[192] = 8'd186;
    sbox_15[193] = 8'd120;
    sbox_15[194] = 8'd37;
    sbox_15[195] = 8'd46;
    sbox_15[196] = 8'd28;
    sbox_15[197] = 8'd166;
    sbox_15[198] = 8'd180;
    sbox_15[199] = 8'd198;
    sbox_15[200] = 8'd232;
    sbox_15[201] = 8'd221;
    sbox_15[202] = 8'd116;
    sbox_15[203] = 8'd31;
    sbox_15[204] = 8'd75;
    sbox_15[205] = 8'd189;
    sbox_15[206] = 8'd139;
    sbox_15[207] = 8'd138;
    sbox_15[208] = 8'd112;
    sbox_15[209] = 8'd62;
    sbox_15[210] = 8'd181;
    sbox_15[211] = 8'd102;
    sbox_15[212] = 8'd72;
    sbox_15[213] = 8'd3;
    sbox_15[214] = 8'd246;
    sbox_15[215] = 8'd14;
    sbox_15[216] = 8'd97;
    sbox_15[217] = 8'd53;
    sbox_15[218] = 8'd87;
    sbox_15[219] = 8'd185;
    sbox_15[220] = 8'd134;
    sbox_15[221] = 8'd193;
    sbox_15[222] = 8'd29;
    sbox_15[223] = 8'd158;
    sbox_15[224] = 8'd225;
    sbox_15[225] = 8'd248;
    sbox_15[226] = 8'd152;
    sbox_15[227] = 8'd17;
    sbox_15[228] = 8'd105;
    sbox_15[229] = 8'd217;
    sbox_15[230] = 8'd142;
    sbox_15[231] = 8'd148;
    sbox_15[232] = 8'd155;
    sbox_15[233] = 8'd30;
    sbox_15[234] = 8'd135;
    sbox_15[235] = 8'd233;
    sbox_15[236] = 8'd206;
    sbox_15[237] = 8'd85;
    sbox_15[238] = 8'd40;
    sbox_15[239] = 8'd223;
    sbox_15[240] = 8'd140;
    sbox_15[241] = 8'd161;
    sbox_15[242] = 8'd137;
    sbox_15[243] = 8'd13;
    sbox_15[244] = 8'd191;
    sbox_15[245] = 8'd230;
    sbox_15[246] = 8'd66;
    sbox_15[247] = 8'd104;
    sbox_15[248] = 8'd65;
    sbox_15[249] = 8'd153;
    sbox_15[250] = 8'd45;
    sbox_15[251] = 8'd15;
    sbox_15[252] = 8'd176;
    sbox_15[253] = 8'd84;
    sbox_15[254] = 8'd187;
    sbox_15[255] = 8'd22;
    sbox_16[0] = 8'd99;
    sbox_16[1] = 8'd124;
    sbox_16[2] = 8'd119;
    sbox_16[3] = 8'd123;
    sbox_16[4] = 8'd242;
    sbox_16[5] = 8'd107;
    sbox_16[6] = 8'd111;
    sbox_16[7] = 8'd197;
    sbox_16[8] = 8'd48;
    sbox_16[9] = 8'd1;
    sbox_16[10] = 8'd103;
    sbox_16[11] = 8'd43;
    sbox_16[12] = 8'd254;
    sbox_16[13] = 8'd215;
    sbox_16[14] = 8'd171;
    sbox_16[15] = 8'd118;
    sbox_16[16] = 8'd202;
    sbox_16[17] = 8'd130;
    sbox_16[18] = 8'd201;
    sbox_16[19] = 8'd125;
    sbox_16[20] = 8'd250;
    sbox_16[21] = 8'd89;
    sbox_16[22] = 8'd71;
    sbox_16[23] = 8'd240;
    sbox_16[24] = 8'd173;
    sbox_16[25] = 8'd212;
    sbox_16[26] = 8'd162;
    sbox_16[27] = 8'd175;
    sbox_16[28] = 8'd156;
    sbox_16[29] = 8'd164;
    sbox_16[30] = 8'd114;
    sbox_16[31] = 8'd192;
    sbox_16[32] = 8'd183;
    sbox_16[33] = 8'd253;
    sbox_16[34] = 8'd147;
    sbox_16[35] = 8'd38;
    sbox_16[36] = 8'd54;
    sbox_16[37] = 8'd63;
    sbox_16[38] = 8'd247;
    sbox_16[39] = 8'd204;
    sbox_16[40] = 8'd52;
    sbox_16[41] = 8'd165;
    sbox_16[42] = 8'd229;
    sbox_16[43] = 8'd241;
    sbox_16[44] = 8'd113;
    sbox_16[45] = 8'd216;
    sbox_16[46] = 8'd49;
    sbox_16[47] = 8'd21;
    sbox_16[48] = 8'd4;
    sbox_16[49] = 8'd199;
    sbox_16[50] = 8'd35;
    sbox_16[51] = 8'd195;
    sbox_16[52] = 8'd24;
    sbox_16[53] = 8'd150;
    sbox_16[54] = 8'd5;
    sbox_16[55] = 8'd154;
    sbox_16[56] = 8'd7;
    sbox_16[57] = 8'd18;
    sbox_16[58] = 8'd128;
    sbox_16[59] = 8'd226;
    sbox_16[60] = 8'd235;
    sbox_16[61] = 8'd39;
    sbox_16[62] = 8'd178;
    sbox_16[63] = 8'd117;
    sbox_16[64] = 8'd9;
    sbox_16[65] = 8'd131;
    sbox_16[66] = 8'd44;
    sbox_16[67] = 8'd26;
    sbox_16[68] = 8'd27;
    sbox_16[69] = 8'd110;
    sbox_16[70] = 8'd90;
    sbox_16[71] = 8'd160;
    sbox_16[72] = 8'd82;
    sbox_16[73] = 8'd59;
    sbox_16[74] = 8'd214;
    sbox_16[75] = 8'd179;
    sbox_16[76] = 8'd41;
    sbox_16[77] = 8'd227;
    sbox_16[78] = 8'd47;
    sbox_16[79] = 8'd132;
    sbox_16[80] = 8'd83;
    sbox_16[81] = 8'd209;
    sbox_16[82] = 8'd0;
    sbox_16[83] = 8'd237;
    sbox_16[84] = 8'd32;
    sbox_16[85] = 8'd252;
    sbox_16[86] = 8'd177;
    sbox_16[87] = 8'd91;
    sbox_16[88] = 8'd106;
    sbox_16[89] = 8'd203;
    sbox_16[90] = 8'd190;
    sbox_16[91] = 8'd57;
    sbox_16[92] = 8'd74;
    sbox_16[93] = 8'd76;
    sbox_16[94] = 8'd88;
    sbox_16[95] = 8'd207;
    sbox_16[96] = 8'd208;
    sbox_16[97] = 8'd239;
    sbox_16[98] = 8'd170;
    sbox_16[99] = 8'd251;
    sbox_16[100] = 8'd67;
    sbox_16[101] = 8'd77;
    sbox_16[102] = 8'd51;
    sbox_16[103] = 8'd133;
    sbox_16[104] = 8'd69;
    sbox_16[105] = 8'd249;
    sbox_16[106] = 8'd2;
    sbox_16[107] = 8'd127;
    sbox_16[108] = 8'd80;
    sbox_16[109] = 8'd60;
    sbox_16[110] = 8'd159;
    sbox_16[111] = 8'd168;
    sbox_16[112] = 8'd81;
    sbox_16[113] = 8'd163;
    sbox_16[114] = 8'd64;
    sbox_16[115] = 8'd143;
    sbox_16[116] = 8'd146;
    sbox_16[117] = 8'd157;
    sbox_16[118] = 8'd56;
    sbox_16[119] = 8'd245;
    sbox_16[120] = 8'd188;
    sbox_16[121] = 8'd182;
    sbox_16[122] = 8'd218;
    sbox_16[123] = 8'd33;
    sbox_16[124] = 8'd16;
    sbox_16[125] = 8'd255;
    sbox_16[126] = 8'd243;
    sbox_16[127] = 8'd210;
    sbox_16[128] = 8'd205;
    sbox_16[129] = 8'd12;
    sbox_16[130] = 8'd19;
    sbox_16[131] = 8'd236;
    sbox_16[132] = 8'd95;
    sbox_16[133] = 8'd151;
    sbox_16[134] = 8'd68;
    sbox_16[135] = 8'd23;
    sbox_16[136] = 8'd196;
    sbox_16[137] = 8'd167;
    sbox_16[138] = 8'd126;
    sbox_16[139] = 8'd61;
    sbox_16[140] = 8'd100;
    sbox_16[141] = 8'd93;
    sbox_16[142] = 8'd25;
    sbox_16[143] = 8'd115;
    sbox_16[144] = 8'd96;
    sbox_16[145] = 8'd129;
    sbox_16[146] = 8'd79;
    sbox_16[147] = 8'd220;
    sbox_16[148] = 8'd34;
    sbox_16[149] = 8'd42;
    sbox_16[150] = 8'd144;
    sbox_16[151] = 8'd136;
    sbox_16[152] = 8'd70;
    sbox_16[153] = 8'd238;
    sbox_16[154] = 8'd184;
    sbox_16[155] = 8'd20;
    sbox_16[156] = 8'd222;
    sbox_16[157] = 8'd94;
    sbox_16[158] = 8'd11;
    sbox_16[159] = 8'd219;
    sbox_16[160] = 8'd224;
    sbox_16[161] = 8'd50;
    sbox_16[162] = 8'd58;
    sbox_16[163] = 8'd10;
    sbox_16[164] = 8'd73;
    sbox_16[165] = 8'd6;
    sbox_16[166] = 8'd36;
    sbox_16[167] = 8'd92;
    sbox_16[168] = 8'd194;
    sbox_16[169] = 8'd211;
    sbox_16[170] = 8'd172;
    sbox_16[171] = 8'd98;
    sbox_16[172] = 8'd145;
    sbox_16[173] = 8'd149;
    sbox_16[174] = 8'd228;
    sbox_16[175] = 8'd121;
    sbox_16[176] = 8'd231;
    sbox_16[177] = 8'd200;
    sbox_16[178] = 8'd55;
    sbox_16[179] = 8'd109;
    sbox_16[180] = 8'd141;
    sbox_16[181] = 8'd213;
    sbox_16[182] = 8'd78;
    sbox_16[183] = 8'd169;
    sbox_16[184] = 8'd108;
    sbox_16[185] = 8'd86;
    sbox_16[186] = 8'd244;
    sbox_16[187] = 8'd234;
    sbox_16[188] = 8'd101;
    sbox_16[189] = 8'd122;
    sbox_16[190] = 8'd174;
    sbox_16[191] = 8'd8;
    sbox_16[192] = 8'd186;
    sbox_16[193] = 8'd120;
    sbox_16[194] = 8'd37;
    sbox_16[195] = 8'd46;
    sbox_16[196] = 8'd28;
    sbox_16[197] = 8'd166;
    sbox_16[198] = 8'd180;
    sbox_16[199] = 8'd198;
    sbox_16[200] = 8'd232;
    sbox_16[201] = 8'd221;
    sbox_16[202] = 8'd116;
    sbox_16[203] = 8'd31;
    sbox_16[204] = 8'd75;
    sbox_16[205] = 8'd189;
    sbox_16[206] = 8'd139;
    sbox_16[207] = 8'd138;
    sbox_16[208] = 8'd112;
    sbox_16[209] = 8'd62;
    sbox_16[210] = 8'd181;
    sbox_16[211] = 8'd102;
    sbox_16[212] = 8'd72;
    sbox_16[213] = 8'd3;
    sbox_16[214] = 8'd246;
    sbox_16[215] = 8'd14;
    sbox_16[216] = 8'd97;
    sbox_16[217] = 8'd53;
    sbox_16[218] = 8'd87;
    sbox_16[219] = 8'd185;
    sbox_16[220] = 8'd134;
    sbox_16[221] = 8'd193;
    sbox_16[222] = 8'd29;
    sbox_16[223] = 8'd158;
    sbox_16[224] = 8'd225;
    sbox_16[225] = 8'd248;
    sbox_16[226] = 8'd152;
    sbox_16[227] = 8'd17;
    sbox_16[228] = 8'd105;
    sbox_16[229] = 8'd217;
    sbox_16[230] = 8'd142;
    sbox_16[231] = 8'd148;
    sbox_16[232] = 8'd155;
    sbox_16[233] = 8'd30;
    sbox_16[234] = 8'd135;
    sbox_16[235] = 8'd233;
    sbox_16[236] = 8'd206;
    sbox_16[237] = 8'd85;
    sbox_16[238] = 8'd40;
    sbox_16[239] = 8'd223;
    sbox_16[240] = 8'd140;
    sbox_16[241] = 8'd161;
    sbox_16[242] = 8'd137;
    sbox_16[243] = 8'd13;
    sbox_16[244] = 8'd191;
    sbox_16[245] = 8'd230;
    sbox_16[246] = 8'd66;
    sbox_16[247] = 8'd104;
    sbox_16[248] = 8'd65;
    sbox_16[249] = 8'd153;
    sbox_16[250] = 8'd45;
    sbox_16[251] = 8'd15;
    sbox_16[252] = 8'd176;
    sbox_16[253] = 8'd84;
    sbox_16[254] = 8'd187;
    sbox_16[255] = 8'd22;
    sbox_17[0] = 8'd99;
    sbox_17[1] = 8'd124;
    sbox_17[2] = 8'd119;
    sbox_17[3] = 8'd123;
    sbox_17[4] = 8'd242;
    sbox_17[5] = 8'd107;
    sbox_17[6] = 8'd111;
    sbox_17[7] = 8'd197;
    sbox_17[8] = 8'd48;
    sbox_17[9] = 8'd1;
    sbox_17[10] = 8'd103;
    sbox_17[11] = 8'd43;
    sbox_17[12] = 8'd254;
    sbox_17[13] = 8'd215;
    sbox_17[14] = 8'd171;
    sbox_17[15] = 8'd118;
    sbox_17[16] = 8'd202;
    sbox_17[17] = 8'd130;
    sbox_17[18] = 8'd201;
    sbox_17[19] = 8'd125;
    sbox_17[20] = 8'd250;
    sbox_17[21] = 8'd89;
    sbox_17[22] = 8'd71;
    sbox_17[23] = 8'd240;
    sbox_17[24] = 8'd173;
    sbox_17[25] = 8'd212;
    sbox_17[26] = 8'd162;
    sbox_17[27] = 8'd175;
    sbox_17[28] = 8'd156;
    sbox_17[29] = 8'd164;
    sbox_17[30] = 8'd114;
    sbox_17[31] = 8'd192;
    sbox_17[32] = 8'd183;
    sbox_17[33] = 8'd253;
    sbox_17[34] = 8'd147;
    sbox_17[35] = 8'd38;
    sbox_17[36] = 8'd54;
    sbox_17[37] = 8'd63;
    sbox_17[38] = 8'd247;
    sbox_17[39] = 8'd204;
    sbox_17[40] = 8'd52;
    sbox_17[41] = 8'd165;
    sbox_17[42] = 8'd229;
    sbox_17[43] = 8'd241;
    sbox_17[44] = 8'd113;
    sbox_17[45] = 8'd216;
    sbox_17[46] = 8'd49;
    sbox_17[47] = 8'd21;
    sbox_17[48] = 8'd4;
    sbox_17[49] = 8'd199;
    sbox_17[50] = 8'd35;
    sbox_17[51] = 8'd195;
    sbox_17[52] = 8'd24;
    sbox_17[53] = 8'd150;
    sbox_17[54] = 8'd5;
    sbox_17[55] = 8'd154;
    sbox_17[56] = 8'd7;
    sbox_17[57] = 8'd18;
    sbox_17[58] = 8'd128;
    sbox_17[59] = 8'd226;
    sbox_17[60] = 8'd235;
    sbox_17[61] = 8'd39;
    sbox_17[62] = 8'd178;
    sbox_17[63] = 8'd117;
    sbox_17[64] = 8'd9;
    sbox_17[65] = 8'd131;
    sbox_17[66] = 8'd44;
    sbox_17[67] = 8'd26;
    sbox_17[68] = 8'd27;
    sbox_17[69] = 8'd110;
    sbox_17[70] = 8'd90;
    sbox_17[71] = 8'd160;
    sbox_17[72] = 8'd82;
    sbox_17[73] = 8'd59;
    sbox_17[74] = 8'd214;
    sbox_17[75] = 8'd179;
    sbox_17[76] = 8'd41;
    sbox_17[77] = 8'd227;
    sbox_17[78] = 8'd47;
    sbox_17[79] = 8'd132;
    sbox_17[80] = 8'd83;
    sbox_17[81] = 8'd209;
    sbox_17[82] = 8'd0;
    sbox_17[83] = 8'd237;
    sbox_17[84] = 8'd32;
    sbox_17[85] = 8'd252;
    sbox_17[86] = 8'd177;
    sbox_17[87] = 8'd91;
    sbox_17[88] = 8'd106;
    sbox_17[89] = 8'd203;
    sbox_17[90] = 8'd190;
    sbox_17[91] = 8'd57;
    sbox_17[92] = 8'd74;
    sbox_17[93] = 8'd76;
    sbox_17[94] = 8'd88;
    sbox_17[95] = 8'd207;
    sbox_17[96] = 8'd208;
    sbox_17[97] = 8'd239;
    sbox_17[98] = 8'd170;
    sbox_17[99] = 8'd251;
    sbox_17[100] = 8'd67;
    sbox_17[101] = 8'd77;
    sbox_17[102] = 8'd51;
    sbox_17[103] = 8'd133;
    sbox_17[104] = 8'd69;
    sbox_17[105] = 8'd249;
    sbox_17[106] = 8'd2;
    sbox_17[107] = 8'd127;
    sbox_17[108] = 8'd80;
    sbox_17[109] = 8'd60;
    sbox_17[110] = 8'd159;
    sbox_17[111] = 8'd168;
    sbox_17[112] = 8'd81;
    sbox_17[113] = 8'd163;
    sbox_17[114] = 8'd64;
    sbox_17[115] = 8'd143;
    sbox_17[116] = 8'd146;
    sbox_17[117] = 8'd157;
    sbox_17[118] = 8'd56;
    sbox_17[119] = 8'd245;
    sbox_17[120] = 8'd188;
    sbox_17[121] = 8'd182;
    sbox_17[122] = 8'd218;
    sbox_17[123] = 8'd33;
    sbox_17[124] = 8'd16;
    sbox_17[125] = 8'd255;
    sbox_17[126] = 8'd243;
    sbox_17[127] = 8'd210;
    sbox_17[128] = 8'd205;
    sbox_17[129] = 8'd12;
    sbox_17[130] = 8'd19;
    sbox_17[131] = 8'd236;
    sbox_17[132] = 8'd95;
    sbox_17[133] = 8'd151;
    sbox_17[134] = 8'd68;
    sbox_17[135] = 8'd23;
    sbox_17[136] = 8'd196;
    sbox_17[137] = 8'd167;
    sbox_17[138] = 8'd126;
    sbox_17[139] = 8'd61;
    sbox_17[140] = 8'd100;
    sbox_17[141] = 8'd93;
    sbox_17[142] = 8'd25;
    sbox_17[143] = 8'd115;
    sbox_17[144] = 8'd96;
    sbox_17[145] = 8'd129;
    sbox_17[146] = 8'd79;
    sbox_17[147] = 8'd220;
    sbox_17[148] = 8'd34;
    sbox_17[149] = 8'd42;
    sbox_17[150] = 8'd144;
    sbox_17[151] = 8'd136;
    sbox_17[152] = 8'd70;
    sbox_17[153] = 8'd238;
    sbox_17[154] = 8'd184;
    sbox_17[155] = 8'd20;
    sbox_17[156] = 8'd222;
    sbox_17[157] = 8'd94;
    sbox_17[158] = 8'd11;
    sbox_17[159] = 8'd219;
    sbox_17[160] = 8'd224;
    sbox_17[161] = 8'd50;
    sbox_17[162] = 8'd58;
    sbox_17[163] = 8'd10;
    sbox_17[164] = 8'd73;
    sbox_17[165] = 8'd6;
    sbox_17[166] = 8'd36;
    sbox_17[167] = 8'd92;
    sbox_17[168] = 8'd194;
    sbox_17[169] = 8'd211;
    sbox_17[170] = 8'd172;
    sbox_17[171] = 8'd98;
    sbox_17[172] = 8'd145;
    sbox_17[173] = 8'd149;
    sbox_17[174] = 8'd228;
    sbox_17[175] = 8'd121;
    sbox_17[176] = 8'd231;
    sbox_17[177] = 8'd200;
    sbox_17[178] = 8'd55;
    sbox_17[179] = 8'd109;
    sbox_17[180] = 8'd141;
    sbox_17[181] = 8'd213;
    sbox_17[182] = 8'd78;
    sbox_17[183] = 8'd169;
    sbox_17[184] = 8'd108;
    sbox_17[185] = 8'd86;
    sbox_17[186] = 8'd244;
    sbox_17[187] = 8'd234;
    sbox_17[188] = 8'd101;
    sbox_17[189] = 8'd122;
    sbox_17[190] = 8'd174;
    sbox_17[191] = 8'd8;
    sbox_17[192] = 8'd186;
    sbox_17[193] = 8'd120;
    sbox_17[194] = 8'd37;
    sbox_17[195] = 8'd46;
    sbox_17[196] = 8'd28;
    sbox_17[197] = 8'd166;
    sbox_17[198] = 8'd180;
    sbox_17[199] = 8'd198;
    sbox_17[200] = 8'd232;
    sbox_17[201] = 8'd221;
    sbox_17[202] = 8'd116;
    sbox_17[203] = 8'd31;
    sbox_17[204] = 8'd75;
    sbox_17[205] = 8'd189;
    sbox_17[206] = 8'd139;
    sbox_17[207] = 8'd138;
    sbox_17[208] = 8'd112;
    sbox_17[209] = 8'd62;
    sbox_17[210] = 8'd181;
    sbox_17[211] = 8'd102;
    sbox_17[212] = 8'd72;
    sbox_17[213] = 8'd3;
    sbox_17[214] = 8'd246;
    sbox_17[215] = 8'd14;
    sbox_17[216] = 8'd97;
    sbox_17[217] = 8'd53;
    sbox_17[218] = 8'd87;
    sbox_17[219] = 8'd185;
    sbox_17[220] = 8'd134;
    sbox_17[221] = 8'd193;
    sbox_17[222] = 8'd29;
    sbox_17[223] = 8'd158;
    sbox_17[224] = 8'd225;
    sbox_17[225] = 8'd248;
    sbox_17[226] = 8'd152;
    sbox_17[227] = 8'd17;
    sbox_17[228] = 8'd105;
    sbox_17[229] = 8'd217;
    sbox_17[230] = 8'd142;
    sbox_17[231] = 8'd148;
    sbox_17[232] = 8'd155;
    sbox_17[233] = 8'd30;
    sbox_17[234] = 8'd135;
    sbox_17[235] = 8'd233;
    sbox_17[236] = 8'd206;
    sbox_17[237] = 8'd85;
    sbox_17[238] = 8'd40;
    sbox_17[239] = 8'd223;
    sbox_17[240] = 8'd140;
    sbox_17[241] = 8'd161;
    sbox_17[242] = 8'd137;
    sbox_17[243] = 8'd13;
    sbox_17[244] = 8'd191;
    sbox_17[245] = 8'd230;
    sbox_17[246] = 8'd66;
    sbox_17[247] = 8'd104;
    sbox_17[248] = 8'd65;
    sbox_17[249] = 8'd153;
    sbox_17[250] = 8'd45;
    sbox_17[251] = 8'd15;
    sbox_17[252] = 8'd176;
    sbox_17[253] = 8'd84;
    sbox_17[254] = 8'd187;
    sbox_17[255] = 8'd22;
    sbox_18[0] = 8'd99;
    sbox_18[1] = 8'd124;
    sbox_18[2] = 8'd119;
    sbox_18[3] = 8'd123;
    sbox_18[4] = 8'd242;
    sbox_18[5] = 8'd107;
    sbox_18[6] = 8'd111;
    sbox_18[7] = 8'd197;
    sbox_18[8] = 8'd48;
    sbox_18[9] = 8'd1;
    sbox_18[10] = 8'd103;
    sbox_18[11] = 8'd43;
    sbox_18[12] = 8'd254;
    sbox_18[13] = 8'd215;
    sbox_18[14] = 8'd171;
    sbox_18[15] = 8'd118;
    sbox_18[16] = 8'd202;
    sbox_18[17] = 8'd130;
    sbox_18[18] = 8'd201;
    sbox_18[19] = 8'd125;
    sbox_18[20] = 8'd250;
    sbox_18[21] = 8'd89;
    sbox_18[22] = 8'd71;
    sbox_18[23] = 8'd240;
    sbox_18[24] = 8'd173;
    sbox_18[25] = 8'd212;
    sbox_18[26] = 8'd162;
    sbox_18[27] = 8'd175;
    sbox_18[28] = 8'd156;
    sbox_18[29] = 8'd164;
    sbox_18[30] = 8'd114;
    sbox_18[31] = 8'd192;
    sbox_18[32] = 8'd183;
    sbox_18[33] = 8'd253;
    sbox_18[34] = 8'd147;
    sbox_18[35] = 8'd38;
    sbox_18[36] = 8'd54;
    sbox_18[37] = 8'd63;
    sbox_18[38] = 8'd247;
    sbox_18[39] = 8'd204;
    sbox_18[40] = 8'd52;
    sbox_18[41] = 8'd165;
    sbox_18[42] = 8'd229;
    sbox_18[43] = 8'd241;
    sbox_18[44] = 8'd113;
    sbox_18[45] = 8'd216;
    sbox_18[46] = 8'd49;
    sbox_18[47] = 8'd21;
    sbox_18[48] = 8'd4;
    sbox_18[49] = 8'd199;
    sbox_18[50] = 8'd35;
    sbox_18[51] = 8'd195;
    sbox_18[52] = 8'd24;
    sbox_18[53] = 8'd150;
    sbox_18[54] = 8'd5;
    sbox_18[55] = 8'd154;
    sbox_18[56] = 8'd7;
    sbox_18[57] = 8'd18;
    sbox_18[58] = 8'd128;
    sbox_18[59] = 8'd226;
    sbox_18[60] = 8'd235;
    sbox_18[61] = 8'd39;
    sbox_18[62] = 8'd178;
    sbox_18[63] = 8'd117;
    sbox_18[64] = 8'd9;
    sbox_18[65] = 8'd131;
    sbox_18[66] = 8'd44;
    sbox_18[67] = 8'd26;
    sbox_18[68] = 8'd27;
    sbox_18[69] = 8'd110;
    sbox_18[70] = 8'd90;
    sbox_18[71] = 8'd160;
    sbox_18[72] = 8'd82;
    sbox_18[73] = 8'd59;
    sbox_18[74] = 8'd214;
    sbox_18[75] = 8'd179;
    sbox_18[76] = 8'd41;
    sbox_18[77] = 8'd227;
    sbox_18[78] = 8'd47;
    sbox_18[79] = 8'd132;
    sbox_18[80] = 8'd83;
    sbox_18[81] = 8'd209;
    sbox_18[82] = 8'd0;
    sbox_18[83] = 8'd237;
    sbox_18[84] = 8'd32;
    sbox_18[85] = 8'd252;
    sbox_18[86] = 8'd177;
    sbox_18[87] = 8'd91;
    sbox_18[88] = 8'd106;
    sbox_18[89] = 8'd203;
    sbox_18[90] = 8'd190;
    sbox_18[91] = 8'd57;
    sbox_18[92] = 8'd74;
    sbox_18[93] = 8'd76;
    sbox_18[94] = 8'd88;
    sbox_18[95] = 8'd207;
    sbox_18[96] = 8'd208;
    sbox_18[97] = 8'd239;
    sbox_18[98] = 8'd170;
    sbox_18[99] = 8'd251;
    sbox_18[100] = 8'd67;
    sbox_18[101] = 8'd77;
    sbox_18[102] = 8'd51;
    sbox_18[103] = 8'd133;
    sbox_18[104] = 8'd69;
    sbox_18[105] = 8'd249;
    sbox_18[106] = 8'd2;
    sbox_18[107] = 8'd127;
    sbox_18[108] = 8'd80;
    sbox_18[109] = 8'd60;
    sbox_18[110] = 8'd159;
    sbox_18[111] = 8'd168;
    sbox_18[112] = 8'd81;
    sbox_18[113] = 8'd163;
    sbox_18[114] = 8'd64;
    sbox_18[115] = 8'd143;
    sbox_18[116] = 8'd146;
    sbox_18[117] = 8'd157;
    sbox_18[118] = 8'd56;
    sbox_18[119] = 8'd245;
    sbox_18[120] = 8'd188;
    sbox_18[121] = 8'd182;
    sbox_18[122] = 8'd218;
    sbox_18[123] = 8'd33;
    sbox_18[124] = 8'd16;
    sbox_18[125] = 8'd255;
    sbox_18[126] = 8'd243;
    sbox_18[127] = 8'd210;
    sbox_18[128] = 8'd205;
    sbox_18[129] = 8'd12;
    sbox_18[130] = 8'd19;
    sbox_18[131] = 8'd236;
    sbox_18[132] = 8'd95;
    sbox_18[133] = 8'd151;
    sbox_18[134] = 8'd68;
    sbox_18[135] = 8'd23;
    sbox_18[136] = 8'd196;
    sbox_18[137] = 8'd167;
    sbox_18[138] = 8'd126;
    sbox_18[139] = 8'd61;
    sbox_18[140] = 8'd100;
    sbox_18[141] = 8'd93;
    sbox_18[142] = 8'd25;
    sbox_18[143] = 8'd115;
    sbox_18[144] = 8'd96;
    sbox_18[145] = 8'd129;
    sbox_18[146] = 8'd79;
    sbox_18[147] = 8'd220;
    sbox_18[148] = 8'd34;
    sbox_18[149] = 8'd42;
    sbox_18[150] = 8'd144;
    sbox_18[151] = 8'd136;
    sbox_18[152] = 8'd70;
    sbox_18[153] = 8'd238;
    sbox_18[154] = 8'd184;
    sbox_18[155] = 8'd20;
    sbox_18[156] = 8'd222;
    sbox_18[157] = 8'd94;
    sbox_18[158] = 8'd11;
    sbox_18[159] = 8'd219;
    sbox_18[160] = 8'd224;
    sbox_18[161] = 8'd50;
    sbox_18[162] = 8'd58;
    sbox_18[163] = 8'd10;
    sbox_18[164] = 8'd73;
    sbox_18[165] = 8'd6;
    sbox_18[166] = 8'd36;
    sbox_18[167] = 8'd92;
    sbox_18[168] = 8'd194;
    sbox_18[169] = 8'd211;
    sbox_18[170] = 8'd172;
    sbox_18[171] = 8'd98;
    sbox_18[172] = 8'd145;
    sbox_18[173] = 8'd149;
    sbox_18[174] = 8'd228;
    sbox_18[175] = 8'd121;
    sbox_18[176] = 8'd231;
    sbox_18[177] = 8'd200;
    sbox_18[178] = 8'd55;
    sbox_18[179] = 8'd109;
    sbox_18[180] = 8'd141;
    sbox_18[181] = 8'd213;
    sbox_18[182] = 8'd78;
    sbox_18[183] = 8'd169;
    sbox_18[184] = 8'd108;
    sbox_18[185] = 8'd86;
    sbox_18[186] = 8'd244;
    sbox_18[187] = 8'd234;
    sbox_18[188] = 8'd101;
    sbox_18[189] = 8'd122;
    sbox_18[190] = 8'd174;
    sbox_18[191] = 8'd8;
    sbox_18[192] = 8'd186;
    sbox_18[193] = 8'd120;
    sbox_18[194] = 8'd37;
    sbox_18[195] = 8'd46;
    sbox_18[196] = 8'd28;
    sbox_18[197] = 8'd166;
    sbox_18[198] = 8'd180;
    sbox_18[199] = 8'd198;
    sbox_18[200] = 8'd232;
    sbox_18[201] = 8'd221;
    sbox_18[202] = 8'd116;
    sbox_18[203] = 8'd31;
    sbox_18[204] = 8'd75;
    sbox_18[205] = 8'd189;
    sbox_18[206] = 8'd139;
    sbox_18[207] = 8'd138;
    sbox_18[208] = 8'd112;
    sbox_18[209] = 8'd62;
    sbox_18[210] = 8'd181;
    sbox_18[211] = 8'd102;
    sbox_18[212] = 8'd72;
    sbox_18[213] = 8'd3;
    sbox_18[214] = 8'd246;
    sbox_18[215] = 8'd14;
    sbox_18[216] = 8'd97;
    sbox_18[217] = 8'd53;
    sbox_18[218] = 8'd87;
    sbox_18[219] = 8'd185;
    sbox_18[220] = 8'd134;
    sbox_18[221] = 8'd193;
    sbox_18[222] = 8'd29;
    sbox_18[223] = 8'd158;
    sbox_18[224] = 8'd225;
    sbox_18[225] = 8'd248;
    sbox_18[226] = 8'd152;
    sbox_18[227] = 8'd17;
    sbox_18[228] = 8'd105;
    sbox_18[229] = 8'd217;
    sbox_18[230] = 8'd142;
    sbox_18[231] = 8'd148;
    sbox_18[232] = 8'd155;
    sbox_18[233] = 8'd30;
    sbox_18[234] = 8'd135;
    sbox_18[235] = 8'd233;
    sbox_18[236] = 8'd206;
    sbox_18[237] = 8'd85;
    sbox_18[238] = 8'd40;
    sbox_18[239] = 8'd223;
    sbox_18[240] = 8'd140;
    sbox_18[241] = 8'd161;
    sbox_18[242] = 8'd137;
    sbox_18[243] = 8'd13;
    sbox_18[244] = 8'd191;
    sbox_18[245] = 8'd230;
    sbox_18[246] = 8'd66;
    sbox_18[247] = 8'd104;
    sbox_18[248] = 8'd65;
    sbox_18[249] = 8'd153;
    sbox_18[250] = 8'd45;
    sbox_18[251] = 8'd15;
    sbox_18[252] = 8'd176;
    sbox_18[253] = 8'd84;
    sbox_18[254] = 8'd187;
    sbox_18[255] = 8'd22;
    sbox_19[0] = 8'd99;
    sbox_19[1] = 8'd124;
    sbox_19[2] = 8'd119;
    sbox_19[3] = 8'd123;
    sbox_19[4] = 8'd242;
    sbox_19[5] = 8'd107;
    sbox_19[6] = 8'd111;
    sbox_19[7] = 8'd197;
    sbox_19[8] = 8'd48;
    sbox_19[9] = 8'd1;
    sbox_19[10] = 8'd103;
    sbox_19[11] = 8'd43;
    sbox_19[12] = 8'd254;
    sbox_19[13] = 8'd215;
    sbox_19[14] = 8'd171;
    sbox_19[15] = 8'd118;
    sbox_19[16] = 8'd202;
    sbox_19[17] = 8'd130;
    sbox_19[18] = 8'd201;
    sbox_19[19] = 8'd125;
    sbox_19[20] = 8'd250;
    sbox_19[21] = 8'd89;
    sbox_19[22] = 8'd71;
    sbox_19[23] = 8'd240;
    sbox_19[24] = 8'd173;
    sbox_19[25] = 8'd212;
    sbox_19[26] = 8'd162;
    sbox_19[27] = 8'd175;
    sbox_19[28] = 8'd156;
    sbox_19[29] = 8'd164;
    sbox_19[30] = 8'd114;
    sbox_19[31] = 8'd192;
    sbox_19[32] = 8'd183;
    sbox_19[33] = 8'd253;
    sbox_19[34] = 8'd147;
    sbox_19[35] = 8'd38;
    sbox_19[36] = 8'd54;
    sbox_19[37] = 8'd63;
    sbox_19[38] = 8'd247;
    sbox_19[39] = 8'd204;
    sbox_19[40] = 8'd52;
    sbox_19[41] = 8'd165;
    sbox_19[42] = 8'd229;
    sbox_19[43] = 8'd241;
    sbox_19[44] = 8'd113;
    sbox_19[45] = 8'd216;
    sbox_19[46] = 8'd49;
    sbox_19[47] = 8'd21;
    sbox_19[48] = 8'd4;
    sbox_19[49] = 8'd199;
    sbox_19[50] = 8'd35;
    sbox_19[51] = 8'd195;
    sbox_19[52] = 8'd24;
    sbox_19[53] = 8'd150;
    sbox_19[54] = 8'd5;
    sbox_19[55] = 8'd154;
    sbox_19[56] = 8'd7;
    sbox_19[57] = 8'd18;
    sbox_19[58] = 8'd128;
    sbox_19[59] = 8'd226;
    sbox_19[60] = 8'd235;
    sbox_19[61] = 8'd39;
    sbox_19[62] = 8'd178;
    sbox_19[63] = 8'd117;
    sbox_19[64] = 8'd9;
    sbox_19[65] = 8'd131;
    sbox_19[66] = 8'd44;
    sbox_19[67] = 8'd26;
    sbox_19[68] = 8'd27;
    sbox_19[69] = 8'd110;
    sbox_19[70] = 8'd90;
    sbox_19[71] = 8'd160;
    sbox_19[72] = 8'd82;
    sbox_19[73] = 8'd59;
    sbox_19[74] = 8'd214;
    sbox_19[75] = 8'd179;
    sbox_19[76] = 8'd41;
    sbox_19[77] = 8'd227;
    sbox_19[78] = 8'd47;
    sbox_19[79] = 8'd132;
    sbox_19[80] = 8'd83;
    sbox_19[81] = 8'd209;
    sbox_19[82] = 8'd0;
    sbox_19[83] = 8'd237;
    sbox_19[84] = 8'd32;
    sbox_19[85] = 8'd252;
    sbox_19[86] = 8'd177;
    sbox_19[87] = 8'd91;
    sbox_19[88] = 8'd106;
    sbox_19[89] = 8'd203;
    sbox_19[90] = 8'd190;
    sbox_19[91] = 8'd57;
    sbox_19[92] = 8'd74;
    sbox_19[93] = 8'd76;
    sbox_19[94] = 8'd88;
    sbox_19[95] = 8'd207;
    sbox_19[96] = 8'd208;
    sbox_19[97] = 8'd239;
    sbox_19[98] = 8'd170;
    sbox_19[99] = 8'd251;
    sbox_19[100] = 8'd67;
    sbox_19[101] = 8'd77;
    sbox_19[102] = 8'd51;
    sbox_19[103] = 8'd133;
    sbox_19[104] = 8'd69;
    sbox_19[105] = 8'd249;
    sbox_19[106] = 8'd2;
    sbox_19[107] = 8'd127;
    sbox_19[108] = 8'd80;
    sbox_19[109] = 8'd60;
    sbox_19[110] = 8'd159;
    sbox_19[111] = 8'd168;
    sbox_19[112] = 8'd81;
    sbox_19[113] = 8'd163;
    sbox_19[114] = 8'd64;
    sbox_19[115] = 8'd143;
    sbox_19[116] = 8'd146;
    sbox_19[117] = 8'd157;
    sbox_19[118] = 8'd56;
    sbox_19[119] = 8'd245;
    sbox_19[120] = 8'd188;
    sbox_19[121] = 8'd182;
    sbox_19[122] = 8'd218;
    sbox_19[123] = 8'd33;
    sbox_19[124] = 8'd16;
    sbox_19[125] = 8'd255;
    sbox_19[126] = 8'd243;
    sbox_19[127] = 8'd210;
    sbox_19[128] = 8'd205;
    sbox_19[129] = 8'd12;
    sbox_19[130] = 8'd19;
    sbox_19[131] = 8'd236;
    sbox_19[132] = 8'd95;
    sbox_19[133] = 8'd151;
    sbox_19[134] = 8'd68;
    sbox_19[135] = 8'd23;
    sbox_19[136] = 8'd196;
    sbox_19[137] = 8'd167;
    sbox_19[138] = 8'd126;
    sbox_19[139] = 8'd61;
    sbox_19[140] = 8'd100;
    sbox_19[141] = 8'd93;
    sbox_19[142] = 8'd25;
    sbox_19[143] = 8'd115;
    sbox_19[144] = 8'd96;
    sbox_19[145] = 8'd129;
    sbox_19[146] = 8'd79;
    sbox_19[147] = 8'd220;
    sbox_19[148] = 8'd34;
    sbox_19[149] = 8'd42;
    sbox_19[150] = 8'd144;
    sbox_19[151] = 8'd136;
    sbox_19[152] = 8'd70;
    sbox_19[153] = 8'd238;
    sbox_19[154] = 8'd184;
    sbox_19[155] = 8'd20;
    sbox_19[156] = 8'd222;
    sbox_19[157] = 8'd94;
    sbox_19[158] = 8'd11;
    sbox_19[159] = 8'd219;
    sbox_19[160] = 8'd224;
    sbox_19[161] = 8'd50;
    sbox_19[162] = 8'd58;
    sbox_19[163] = 8'd10;
    sbox_19[164] = 8'd73;
    sbox_19[165] = 8'd6;
    sbox_19[166] = 8'd36;
    sbox_19[167] = 8'd92;
    sbox_19[168] = 8'd194;
    sbox_19[169] = 8'd211;
    sbox_19[170] = 8'd172;
    sbox_19[171] = 8'd98;
    sbox_19[172] = 8'd145;
    sbox_19[173] = 8'd149;
    sbox_19[174] = 8'd228;
    sbox_19[175] = 8'd121;
    sbox_19[176] = 8'd231;
    sbox_19[177] = 8'd200;
    sbox_19[178] = 8'd55;
    sbox_19[179] = 8'd109;
    sbox_19[180] = 8'd141;
    sbox_19[181] = 8'd213;
    sbox_19[182] = 8'd78;
    sbox_19[183] = 8'd169;
    sbox_19[184] = 8'd108;
    sbox_19[185] = 8'd86;
    sbox_19[186] = 8'd244;
    sbox_19[187] = 8'd234;
    sbox_19[188] = 8'd101;
    sbox_19[189] = 8'd122;
    sbox_19[190] = 8'd174;
    sbox_19[191] = 8'd8;
    sbox_19[192] = 8'd186;
    sbox_19[193] = 8'd120;
    sbox_19[194] = 8'd37;
    sbox_19[195] = 8'd46;
    sbox_19[196] = 8'd28;
    sbox_19[197] = 8'd166;
    sbox_19[198] = 8'd180;
    sbox_19[199] = 8'd198;
    sbox_19[200] = 8'd232;
    sbox_19[201] = 8'd221;
    sbox_19[202] = 8'd116;
    sbox_19[203] = 8'd31;
    sbox_19[204] = 8'd75;
    sbox_19[205] = 8'd189;
    sbox_19[206] = 8'd139;
    sbox_19[207] = 8'd138;
    sbox_19[208] = 8'd112;
    sbox_19[209] = 8'd62;
    sbox_19[210] = 8'd181;
    sbox_19[211] = 8'd102;
    sbox_19[212] = 8'd72;
    sbox_19[213] = 8'd3;
    sbox_19[214] = 8'd246;
    sbox_19[215] = 8'd14;
    sbox_19[216] = 8'd97;
    sbox_19[217] = 8'd53;
    sbox_19[218] = 8'd87;
    sbox_19[219] = 8'd185;
    sbox_19[220] = 8'd134;
    sbox_19[221] = 8'd193;
    sbox_19[222] = 8'd29;
    sbox_19[223] = 8'd158;
    sbox_19[224] = 8'd225;
    sbox_19[225] = 8'd248;
    sbox_19[226] = 8'd152;
    sbox_19[227] = 8'd17;
    sbox_19[228] = 8'd105;
    sbox_19[229] = 8'd217;
    sbox_19[230] = 8'd142;
    sbox_19[231] = 8'd148;
    sbox_19[232] = 8'd155;
    sbox_19[233] = 8'd30;
    sbox_19[234] = 8'd135;
    sbox_19[235] = 8'd233;
    sbox_19[236] = 8'd206;
    sbox_19[237] = 8'd85;
    sbox_19[238] = 8'd40;
    sbox_19[239] = 8'd223;
    sbox_19[240] = 8'd140;
    sbox_19[241] = 8'd161;
    sbox_19[242] = 8'd137;
    sbox_19[243] = 8'd13;
    sbox_19[244] = 8'd191;
    sbox_19[245] = 8'd230;
    sbox_19[246] = 8'd66;
    sbox_19[247] = 8'd104;
    sbox_19[248] = 8'd65;
    sbox_19[249] = 8'd153;
    sbox_19[250] = 8'd45;
    sbox_19[251] = 8'd15;
    sbox_19[252] = 8'd176;
    sbox_19[253] = 8'd84;
    sbox_19[254] = 8'd187;
    sbox_19[255] = 8'd22;
    sbox_20[0] = 8'd99;
    sbox_20[1] = 8'd124;
    sbox_20[2] = 8'd119;
    sbox_20[3] = 8'd123;
    sbox_20[4] = 8'd242;
    sbox_20[5] = 8'd107;
    sbox_20[6] = 8'd111;
    sbox_20[7] = 8'd197;
    sbox_20[8] = 8'd48;
    sbox_20[9] = 8'd1;
    sbox_20[10] = 8'd103;
    sbox_20[11] = 8'd43;
    sbox_20[12] = 8'd254;
    sbox_20[13] = 8'd215;
    sbox_20[14] = 8'd171;
    sbox_20[15] = 8'd118;
    sbox_20[16] = 8'd202;
    sbox_20[17] = 8'd130;
    sbox_20[18] = 8'd201;
    sbox_20[19] = 8'd125;
    sbox_20[20] = 8'd250;
    sbox_20[21] = 8'd89;
    sbox_20[22] = 8'd71;
    sbox_20[23] = 8'd240;
    sbox_20[24] = 8'd173;
    sbox_20[25] = 8'd212;
    sbox_20[26] = 8'd162;
    sbox_20[27] = 8'd175;
    sbox_20[28] = 8'd156;
    sbox_20[29] = 8'd164;
    sbox_20[30] = 8'd114;
    sbox_20[31] = 8'd192;
    sbox_20[32] = 8'd183;
    sbox_20[33] = 8'd253;
    sbox_20[34] = 8'd147;
    sbox_20[35] = 8'd38;
    sbox_20[36] = 8'd54;
    sbox_20[37] = 8'd63;
    sbox_20[38] = 8'd247;
    sbox_20[39] = 8'd204;
    sbox_20[40] = 8'd52;
    sbox_20[41] = 8'd165;
    sbox_20[42] = 8'd229;
    sbox_20[43] = 8'd241;
    sbox_20[44] = 8'd113;
    sbox_20[45] = 8'd216;
    sbox_20[46] = 8'd49;
    sbox_20[47] = 8'd21;
    sbox_20[48] = 8'd4;
    sbox_20[49] = 8'd199;
    sbox_20[50] = 8'd35;
    sbox_20[51] = 8'd195;
    sbox_20[52] = 8'd24;
    sbox_20[53] = 8'd150;
    sbox_20[54] = 8'd5;
    sbox_20[55] = 8'd154;
    sbox_20[56] = 8'd7;
    sbox_20[57] = 8'd18;
    sbox_20[58] = 8'd128;
    sbox_20[59] = 8'd226;
    sbox_20[60] = 8'd235;
    sbox_20[61] = 8'd39;
    sbox_20[62] = 8'd178;
    sbox_20[63] = 8'd117;
    sbox_20[64] = 8'd9;
    sbox_20[65] = 8'd131;
    sbox_20[66] = 8'd44;
    sbox_20[67] = 8'd26;
    sbox_20[68] = 8'd27;
    sbox_20[69] = 8'd110;
    sbox_20[70] = 8'd90;
    sbox_20[71] = 8'd160;
    sbox_20[72] = 8'd82;
    sbox_20[73] = 8'd59;
    sbox_20[74] = 8'd214;
    sbox_20[75] = 8'd179;
    sbox_20[76] = 8'd41;
    sbox_20[77] = 8'd227;
    sbox_20[78] = 8'd47;
    sbox_20[79] = 8'd132;
    sbox_20[80] = 8'd83;
    sbox_20[81] = 8'd209;
    sbox_20[82] = 8'd0;
    sbox_20[83] = 8'd237;
    sbox_20[84] = 8'd32;
    sbox_20[85] = 8'd252;
    sbox_20[86] = 8'd177;
    sbox_20[87] = 8'd91;
    sbox_20[88] = 8'd106;
    sbox_20[89] = 8'd203;
    sbox_20[90] = 8'd190;
    sbox_20[91] = 8'd57;
    sbox_20[92] = 8'd74;
    sbox_20[93] = 8'd76;
    sbox_20[94] = 8'd88;
    sbox_20[95] = 8'd207;
    sbox_20[96] = 8'd208;
    sbox_20[97] = 8'd239;
    sbox_20[98] = 8'd170;
    sbox_20[99] = 8'd251;
    sbox_20[100] = 8'd67;
    sbox_20[101] = 8'd77;
    sbox_20[102] = 8'd51;
    sbox_20[103] = 8'd133;
    sbox_20[104] = 8'd69;
    sbox_20[105] = 8'd249;
    sbox_20[106] = 8'd2;
    sbox_20[107] = 8'd127;
    sbox_20[108] = 8'd80;
    sbox_20[109] = 8'd60;
    sbox_20[110] = 8'd159;
    sbox_20[111] = 8'd168;
    sbox_20[112] = 8'd81;
    sbox_20[113] = 8'd163;
    sbox_20[114] = 8'd64;
    sbox_20[115] = 8'd143;
    sbox_20[116] = 8'd146;
    sbox_20[117] = 8'd157;
    sbox_20[118] = 8'd56;
    sbox_20[119] = 8'd245;
    sbox_20[120] = 8'd188;
    sbox_20[121] = 8'd182;
    sbox_20[122] = 8'd218;
    sbox_20[123] = 8'd33;
    sbox_20[124] = 8'd16;
    sbox_20[125] = 8'd255;
    sbox_20[126] = 8'd243;
    sbox_20[127] = 8'd210;
    sbox_20[128] = 8'd205;
    sbox_20[129] = 8'd12;
    sbox_20[130] = 8'd19;
    sbox_20[131] = 8'd236;
    sbox_20[132] = 8'd95;
    sbox_20[133] = 8'd151;
    sbox_20[134] = 8'd68;
    sbox_20[135] = 8'd23;
    sbox_20[136] = 8'd196;
    sbox_20[137] = 8'd167;
    sbox_20[138] = 8'd126;
    sbox_20[139] = 8'd61;
    sbox_20[140] = 8'd100;
    sbox_20[141] = 8'd93;
    sbox_20[142] = 8'd25;
    sbox_20[143] = 8'd115;
    sbox_20[144] = 8'd96;
    sbox_20[145] = 8'd129;
    sbox_20[146] = 8'd79;
    sbox_20[147] = 8'd220;
    sbox_20[148] = 8'd34;
    sbox_20[149] = 8'd42;
    sbox_20[150] = 8'd144;
    sbox_20[151] = 8'd136;
    sbox_20[152] = 8'd70;
    sbox_20[153] = 8'd238;
    sbox_20[154] = 8'd184;
    sbox_20[155] = 8'd20;
    sbox_20[156] = 8'd222;
    sbox_20[157] = 8'd94;
    sbox_20[158] = 8'd11;
    sbox_20[159] = 8'd219;
    sbox_20[160] = 8'd224;
    sbox_20[161] = 8'd50;
    sbox_20[162] = 8'd58;
    sbox_20[163] = 8'd10;
    sbox_20[164] = 8'd73;
    sbox_20[165] = 8'd6;
    sbox_20[166] = 8'd36;
    sbox_20[167] = 8'd92;
    sbox_20[168] = 8'd194;
    sbox_20[169] = 8'd211;
    sbox_20[170] = 8'd172;
    sbox_20[171] = 8'd98;
    sbox_20[172] = 8'd145;
    sbox_20[173] = 8'd149;
    sbox_20[174] = 8'd228;
    sbox_20[175] = 8'd121;
    sbox_20[176] = 8'd231;
    sbox_20[177] = 8'd200;
    sbox_20[178] = 8'd55;
    sbox_20[179] = 8'd109;
    sbox_20[180] = 8'd141;
    sbox_20[181] = 8'd213;
    sbox_20[182] = 8'd78;
    sbox_20[183] = 8'd169;
    sbox_20[184] = 8'd108;
    sbox_20[185] = 8'd86;
    sbox_20[186] = 8'd244;
    sbox_20[187] = 8'd234;
    sbox_20[188] = 8'd101;
    sbox_20[189] = 8'd122;
    sbox_20[190] = 8'd174;
    sbox_20[191] = 8'd8;
    sbox_20[192] = 8'd186;
    sbox_20[193] = 8'd120;
    sbox_20[194] = 8'd37;
    sbox_20[195] = 8'd46;
    sbox_20[196] = 8'd28;
    sbox_20[197] = 8'd166;
    sbox_20[198] = 8'd180;
    sbox_20[199] = 8'd198;
    sbox_20[200] = 8'd232;
    sbox_20[201] = 8'd221;
    sbox_20[202] = 8'd116;
    sbox_20[203] = 8'd31;
    sbox_20[204] = 8'd75;
    sbox_20[205] = 8'd189;
    sbox_20[206] = 8'd139;
    sbox_20[207] = 8'd138;
    sbox_20[208] = 8'd112;
    sbox_20[209] = 8'd62;
    sbox_20[210] = 8'd181;
    sbox_20[211] = 8'd102;
    sbox_20[212] = 8'd72;
    sbox_20[213] = 8'd3;
    sbox_20[214] = 8'd246;
    sbox_20[215] = 8'd14;
    sbox_20[216] = 8'd97;
    sbox_20[217] = 8'd53;
    sbox_20[218] = 8'd87;
    sbox_20[219] = 8'd185;
    sbox_20[220] = 8'd134;
    sbox_20[221] = 8'd193;
    sbox_20[222] = 8'd29;
    sbox_20[223] = 8'd158;
    sbox_20[224] = 8'd225;
    sbox_20[225] = 8'd248;
    sbox_20[226] = 8'd152;
    sbox_20[227] = 8'd17;
    sbox_20[228] = 8'd105;
    sbox_20[229] = 8'd217;
    sbox_20[230] = 8'd142;
    sbox_20[231] = 8'd148;
    sbox_20[232] = 8'd155;
    sbox_20[233] = 8'd30;
    sbox_20[234] = 8'd135;
    sbox_20[235] = 8'd233;
    sbox_20[236] = 8'd206;
    sbox_20[237] = 8'd85;
    sbox_20[238] = 8'd40;
    sbox_20[239] = 8'd223;
    sbox_20[240] = 8'd140;
    sbox_20[241] = 8'd161;
    sbox_20[242] = 8'd137;
    sbox_20[243] = 8'd13;
    sbox_20[244] = 8'd191;
    sbox_20[245] = 8'd230;
    sbox_20[246] = 8'd66;
    sbox_20[247] = 8'd104;
    sbox_20[248] = 8'd65;
    sbox_20[249] = 8'd153;
    sbox_20[250] = 8'd45;
    sbox_20[251] = 8'd15;
    sbox_20[252] = 8'd176;
    sbox_20[253] = 8'd84;
    sbox_20[254] = 8'd187;
    sbox_20[255] = 8'd22;
    sbox_21[0] = 8'd99;
    sbox_21[1] = 8'd124;
    sbox_21[2] = 8'd119;
    sbox_21[3] = 8'd123;
    sbox_21[4] = 8'd242;
    sbox_21[5] = 8'd107;
    sbox_21[6] = 8'd111;
    sbox_21[7] = 8'd197;
    sbox_21[8] = 8'd48;
    sbox_21[9] = 8'd1;
    sbox_21[10] = 8'd103;
    sbox_21[11] = 8'd43;
    sbox_21[12] = 8'd254;
    sbox_21[13] = 8'd215;
    sbox_21[14] = 8'd171;
    sbox_21[15] = 8'd118;
    sbox_21[16] = 8'd202;
    sbox_21[17] = 8'd130;
    sbox_21[18] = 8'd201;
    sbox_21[19] = 8'd125;
    sbox_21[20] = 8'd250;
    sbox_21[21] = 8'd89;
    sbox_21[22] = 8'd71;
    sbox_21[23] = 8'd240;
    sbox_21[24] = 8'd173;
    sbox_21[25] = 8'd212;
    sbox_21[26] = 8'd162;
    sbox_21[27] = 8'd175;
    sbox_21[28] = 8'd156;
    sbox_21[29] = 8'd164;
    sbox_21[30] = 8'd114;
    sbox_21[31] = 8'd192;
    sbox_21[32] = 8'd183;
    sbox_21[33] = 8'd253;
    sbox_21[34] = 8'd147;
    sbox_21[35] = 8'd38;
    sbox_21[36] = 8'd54;
    sbox_21[37] = 8'd63;
    sbox_21[38] = 8'd247;
    sbox_21[39] = 8'd204;
    sbox_21[40] = 8'd52;
    sbox_21[41] = 8'd165;
    sbox_21[42] = 8'd229;
    sbox_21[43] = 8'd241;
    sbox_21[44] = 8'd113;
    sbox_21[45] = 8'd216;
    sbox_21[46] = 8'd49;
    sbox_21[47] = 8'd21;
    sbox_21[48] = 8'd4;
    sbox_21[49] = 8'd199;
    sbox_21[50] = 8'd35;
    sbox_21[51] = 8'd195;
    sbox_21[52] = 8'd24;
    sbox_21[53] = 8'd150;
    sbox_21[54] = 8'd5;
    sbox_21[55] = 8'd154;
    sbox_21[56] = 8'd7;
    sbox_21[57] = 8'd18;
    sbox_21[58] = 8'd128;
    sbox_21[59] = 8'd226;
    sbox_21[60] = 8'd235;
    sbox_21[61] = 8'd39;
    sbox_21[62] = 8'd178;
    sbox_21[63] = 8'd117;
    sbox_21[64] = 8'd9;
    sbox_21[65] = 8'd131;
    sbox_21[66] = 8'd44;
    sbox_21[67] = 8'd26;
    sbox_21[68] = 8'd27;
    sbox_21[69] = 8'd110;
    sbox_21[70] = 8'd90;
    sbox_21[71] = 8'd160;
    sbox_21[72] = 8'd82;
    sbox_21[73] = 8'd59;
    sbox_21[74] = 8'd214;
    sbox_21[75] = 8'd179;
    sbox_21[76] = 8'd41;
    sbox_21[77] = 8'd227;
    sbox_21[78] = 8'd47;
    sbox_21[79] = 8'd132;
    sbox_21[80] = 8'd83;
    sbox_21[81] = 8'd209;
    sbox_21[82] = 8'd0;
    sbox_21[83] = 8'd237;
    sbox_21[84] = 8'd32;
    sbox_21[85] = 8'd252;
    sbox_21[86] = 8'd177;
    sbox_21[87] = 8'd91;
    sbox_21[88] = 8'd106;
    sbox_21[89] = 8'd203;
    sbox_21[90] = 8'd190;
    sbox_21[91] = 8'd57;
    sbox_21[92] = 8'd74;
    sbox_21[93] = 8'd76;
    sbox_21[94] = 8'd88;
    sbox_21[95] = 8'd207;
    sbox_21[96] = 8'd208;
    sbox_21[97] = 8'd239;
    sbox_21[98] = 8'd170;
    sbox_21[99] = 8'd251;
    sbox_21[100] = 8'd67;
    sbox_21[101] = 8'd77;
    sbox_21[102] = 8'd51;
    sbox_21[103] = 8'd133;
    sbox_21[104] = 8'd69;
    sbox_21[105] = 8'd249;
    sbox_21[106] = 8'd2;
    sbox_21[107] = 8'd127;
    sbox_21[108] = 8'd80;
    sbox_21[109] = 8'd60;
    sbox_21[110] = 8'd159;
    sbox_21[111] = 8'd168;
    sbox_21[112] = 8'd81;
    sbox_21[113] = 8'd163;
    sbox_21[114] = 8'd64;
    sbox_21[115] = 8'd143;
    sbox_21[116] = 8'd146;
    sbox_21[117] = 8'd157;
    sbox_21[118] = 8'd56;
    sbox_21[119] = 8'd245;
    sbox_21[120] = 8'd188;
    sbox_21[121] = 8'd182;
    sbox_21[122] = 8'd218;
    sbox_21[123] = 8'd33;
    sbox_21[124] = 8'd16;
    sbox_21[125] = 8'd255;
    sbox_21[126] = 8'd243;
    sbox_21[127] = 8'd210;
    sbox_21[128] = 8'd205;
    sbox_21[129] = 8'd12;
    sbox_21[130] = 8'd19;
    sbox_21[131] = 8'd236;
    sbox_21[132] = 8'd95;
    sbox_21[133] = 8'd151;
    sbox_21[134] = 8'd68;
    sbox_21[135] = 8'd23;
    sbox_21[136] = 8'd196;
    sbox_21[137] = 8'd167;
    sbox_21[138] = 8'd126;
    sbox_21[139] = 8'd61;
    sbox_21[140] = 8'd100;
    sbox_21[141] = 8'd93;
    sbox_21[142] = 8'd25;
    sbox_21[143] = 8'd115;
    sbox_21[144] = 8'd96;
    sbox_21[145] = 8'd129;
    sbox_21[146] = 8'd79;
    sbox_21[147] = 8'd220;
    sbox_21[148] = 8'd34;
    sbox_21[149] = 8'd42;
    sbox_21[150] = 8'd144;
    sbox_21[151] = 8'd136;
    sbox_21[152] = 8'd70;
    sbox_21[153] = 8'd238;
    sbox_21[154] = 8'd184;
    sbox_21[155] = 8'd20;
    sbox_21[156] = 8'd222;
    sbox_21[157] = 8'd94;
    sbox_21[158] = 8'd11;
    sbox_21[159] = 8'd219;
    sbox_21[160] = 8'd224;
    sbox_21[161] = 8'd50;
    sbox_21[162] = 8'd58;
    sbox_21[163] = 8'd10;
    sbox_21[164] = 8'd73;
    sbox_21[165] = 8'd6;
    sbox_21[166] = 8'd36;
    sbox_21[167] = 8'd92;
    sbox_21[168] = 8'd194;
    sbox_21[169] = 8'd211;
    sbox_21[170] = 8'd172;
    sbox_21[171] = 8'd98;
    sbox_21[172] = 8'd145;
    sbox_21[173] = 8'd149;
    sbox_21[174] = 8'd228;
    sbox_21[175] = 8'd121;
    sbox_21[176] = 8'd231;
    sbox_21[177] = 8'd200;
    sbox_21[178] = 8'd55;
    sbox_21[179] = 8'd109;
    sbox_21[180] = 8'd141;
    sbox_21[181] = 8'd213;
    sbox_21[182] = 8'd78;
    sbox_21[183] = 8'd169;
    sbox_21[184] = 8'd108;
    sbox_21[185] = 8'd86;
    sbox_21[186] = 8'd244;
    sbox_21[187] = 8'd234;
    sbox_21[188] = 8'd101;
    sbox_21[189] = 8'd122;
    sbox_21[190] = 8'd174;
    sbox_21[191] = 8'd8;
    sbox_21[192] = 8'd186;
    sbox_21[193] = 8'd120;
    sbox_21[194] = 8'd37;
    sbox_21[195] = 8'd46;
    sbox_21[196] = 8'd28;
    sbox_21[197] = 8'd166;
    sbox_21[198] = 8'd180;
    sbox_21[199] = 8'd198;
    sbox_21[200] = 8'd232;
    sbox_21[201] = 8'd221;
    sbox_21[202] = 8'd116;
    sbox_21[203] = 8'd31;
    sbox_21[204] = 8'd75;
    sbox_21[205] = 8'd189;
    sbox_21[206] = 8'd139;
    sbox_21[207] = 8'd138;
    sbox_21[208] = 8'd112;
    sbox_21[209] = 8'd62;
    sbox_21[210] = 8'd181;
    sbox_21[211] = 8'd102;
    sbox_21[212] = 8'd72;
    sbox_21[213] = 8'd3;
    sbox_21[214] = 8'd246;
    sbox_21[215] = 8'd14;
    sbox_21[216] = 8'd97;
    sbox_21[217] = 8'd53;
    sbox_21[218] = 8'd87;
    sbox_21[219] = 8'd185;
    sbox_21[220] = 8'd134;
    sbox_21[221] = 8'd193;
    sbox_21[222] = 8'd29;
    sbox_21[223] = 8'd158;
    sbox_21[224] = 8'd225;
    sbox_21[225] = 8'd248;
    sbox_21[226] = 8'd152;
    sbox_21[227] = 8'd17;
    sbox_21[228] = 8'd105;
    sbox_21[229] = 8'd217;
    sbox_21[230] = 8'd142;
    sbox_21[231] = 8'd148;
    sbox_21[232] = 8'd155;
    sbox_21[233] = 8'd30;
    sbox_21[234] = 8'd135;
    sbox_21[235] = 8'd233;
    sbox_21[236] = 8'd206;
    sbox_21[237] = 8'd85;
    sbox_21[238] = 8'd40;
    sbox_21[239] = 8'd223;
    sbox_21[240] = 8'd140;
    sbox_21[241] = 8'd161;
    sbox_21[242] = 8'd137;
    sbox_21[243] = 8'd13;
    sbox_21[244] = 8'd191;
    sbox_21[245] = 8'd230;
    sbox_21[246] = 8'd66;
    sbox_21[247] = 8'd104;
    sbox_21[248] = 8'd65;
    sbox_21[249] = 8'd153;
    sbox_21[250] = 8'd45;
    sbox_21[251] = 8'd15;
    sbox_21[252] = 8'd176;
    sbox_21[253] = 8'd84;
    sbox_21[254] = 8'd187;
    sbox_21[255] = 8'd22;
    sbox_22[0] = 8'd99;
    sbox_22[1] = 8'd124;
    sbox_22[2] = 8'd119;
    sbox_22[3] = 8'd123;
    sbox_22[4] = 8'd242;
    sbox_22[5] = 8'd107;
    sbox_22[6] = 8'd111;
    sbox_22[7] = 8'd197;
    sbox_22[8] = 8'd48;
    sbox_22[9] = 8'd1;
    sbox_22[10] = 8'd103;
    sbox_22[11] = 8'd43;
    sbox_22[12] = 8'd254;
    sbox_22[13] = 8'd215;
    sbox_22[14] = 8'd171;
    sbox_22[15] = 8'd118;
    sbox_22[16] = 8'd202;
    sbox_22[17] = 8'd130;
    sbox_22[18] = 8'd201;
    sbox_22[19] = 8'd125;
    sbox_22[20] = 8'd250;
    sbox_22[21] = 8'd89;
    sbox_22[22] = 8'd71;
    sbox_22[23] = 8'd240;
    sbox_22[24] = 8'd173;
    sbox_22[25] = 8'd212;
    sbox_22[26] = 8'd162;
    sbox_22[27] = 8'd175;
    sbox_22[28] = 8'd156;
    sbox_22[29] = 8'd164;
    sbox_22[30] = 8'd114;
    sbox_22[31] = 8'd192;
    sbox_22[32] = 8'd183;
    sbox_22[33] = 8'd253;
    sbox_22[34] = 8'd147;
    sbox_22[35] = 8'd38;
    sbox_22[36] = 8'd54;
    sbox_22[37] = 8'd63;
    sbox_22[38] = 8'd247;
    sbox_22[39] = 8'd204;
    sbox_22[40] = 8'd52;
    sbox_22[41] = 8'd165;
    sbox_22[42] = 8'd229;
    sbox_22[43] = 8'd241;
    sbox_22[44] = 8'd113;
    sbox_22[45] = 8'd216;
    sbox_22[46] = 8'd49;
    sbox_22[47] = 8'd21;
    sbox_22[48] = 8'd4;
    sbox_22[49] = 8'd199;
    sbox_22[50] = 8'd35;
    sbox_22[51] = 8'd195;
    sbox_22[52] = 8'd24;
    sbox_22[53] = 8'd150;
    sbox_22[54] = 8'd5;
    sbox_22[55] = 8'd154;
    sbox_22[56] = 8'd7;
    sbox_22[57] = 8'd18;
    sbox_22[58] = 8'd128;
    sbox_22[59] = 8'd226;
    sbox_22[60] = 8'd235;
    sbox_22[61] = 8'd39;
    sbox_22[62] = 8'd178;
    sbox_22[63] = 8'd117;
    sbox_22[64] = 8'd9;
    sbox_22[65] = 8'd131;
    sbox_22[66] = 8'd44;
    sbox_22[67] = 8'd26;
    sbox_22[68] = 8'd27;
    sbox_22[69] = 8'd110;
    sbox_22[70] = 8'd90;
    sbox_22[71] = 8'd160;
    sbox_22[72] = 8'd82;
    sbox_22[73] = 8'd59;
    sbox_22[74] = 8'd214;
    sbox_22[75] = 8'd179;
    sbox_22[76] = 8'd41;
    sbox_22[77] = 8'd227;
    sbox_22[78] = 8'd47;
    sbox_22[79] = 8'd132;
    sbox_22[80] = 8'd83;
    sbox_22[81] = 8'd209;
    sbox_22[82] = 8'd0;
    sbox_22[83] = 8'd237;
    sbox_22[84] = 8'd32;
    sbox_22[85] = 8'd252;
    sbox_22[86] = 8'd177;
    sbox_22[87] = 8'd91;
    sbox_22[88] = 8'd106;
    sbox_22[89] = 8'd203;
    sbox_22[90] = 8'd190;
    sbox_22[91] = 8'd57;
    sbox_22[92] = 8'd74;
    sbox_22[93] = 8'd76;
    sbox_22[94] = 8'd88;
    sbox_22[95] = 8'd207;
    sbox_22[96] = 8'd208;
    sbox_22[97] = 8'd239;
    sbox_22[98] = 8'd170;
    sbox_22[99] = 8'd251;
    sbox_22[100] = 8'd67;
    sbox_22[101] = 8'd77;
    sbox_22[102] = 8'd51;
    sbox_22[103] = 8'd133;
    sbox_22[104] = 8'd69;
    sbox_22[105] = 8'd249;
    sbox_22[106] = 8'd2;
    sbox_22[107] = 8'd127;
    sbox_22[108] = 8'd80;
    sbox_22[109] = 8'd60;
    sbox_22[110] = 8'd159;
    sbox_22[111] = 8'd168;
    sbox_22[112] = 8'd81;
    sbox_22[113] = 8'd163;
    sbox_22[114] = 8'd64;
    sbox_22[115] = 8'd143;
    sbox_22[116] = 8'd146;
    sbox_22[117] = 8'd157;
    sbox_22[118] = 8'd56;
    sbox_22[119] = 8'd245;
    sbox_22[120] = 8'd188;
    sbox_22[121] = 8'd182;
    sbox_22[122] = 8'd218;
    sbox_22[123] = 8'd33;
    sbox_22[124] = 8'd16;
    sbox_22[125] = 8'd255;
    sbox_22[126] = 8'd243;
    sbox_22[127] = 8'd210;
    sbox_22[128] = 8'd205;
    sbox_22[129] = 8'd12;
    sbox_22[130] = 8'd19;
    sbox_22[131] = 8'd236;
    sbox_22[132] = 8'd95;
    sbox_22[133] = 8'd151;
    sbox_22[134] = 8'd68;
    sbox_22[135] = 8'd23;
    sbox_22[136] = 8'd196;
    sbox_22[137] = 8'd167;
    sbox_22[138] = 8'd126;
    sbox_22[139] = 8'd61;
    sbox_22[140] = 8'd100;
    sbox_22[141] = 8'd93;
    sbox_22[142] = 8'd25;
    sbox_22[143] = 8'd115;
    sbox_22[144] = 8'd96;
    sbox_22[145] = 8'd129;
    sbox_22[146] = 8'd79;
    sbox_22[147] = 8'd220;
    sbox_22[148] = 8'd34;
    sbox_22[149] = 8'd42;
    sbox_22[150] = 8'd144;
    sbox_22[151] = 8'd136;
    sbox_22[152] = 8'd70;
    sbox_22[153] = 8'd238;
    sbox_22[154] = 8'd184;
    sbox_22[155] = 8'd20;
    sbox_22[156] = 8'd222;
    sbox_22[157] = 8'd94;
    sbox_22[158] = 8'd11;
    sbox_22[159] = 8'd219;
    sbox_22[160] = 8'd224;
    sbox_22[161] = 8'd50;
    sbox_22[162] = 8'd58;
    sbox_22[163] = 8'd10;
    sbox_22[164] = 8'd73;
    sbox_22[165] = 8'd6;
    sbox_22[166] = 8'd36;
    sbox_22[167] = 8'd92;
    sbox_22[168] = 8'd194;
    sbox_22[169] = 8'd211;
    sbox_22[170] = 8'd172;
    sbox_22[171] = 8'd98;
    sbox_22[172] = 8'd145;
    sbox_22[173] = 8'd149;
    sbox_22[174] = 8'd228;
    sbox_22[175] = 8'd121;
    sbox_22[176] = 8'd231;
    sbox_22[177] = 8'd200;
    sbox_22[178] = 8'd55;
    sbox_22[179] = 8'd109;
    sbox_22[180] = 8'd141;
    sbox_22[181] = 8'd213;
    sbox_22[182] = 8'd78;
    sbox_22[183] = 8'd169;
    sbox_22[184] = 8'd108;
    sbox_22[185] = 8'd86;
    sbox_22[186] = 8'd244;
    sbox_22[187] = 8'd234;
    sbox_22[188] = 8'd101;
    sbox_22[189] = 8'd122;
    sbox_22[190] = 8'd174;
    sbox_22[191] = 8'd8;
    sbox_22[192] = 8'd186;
    sbox_22[193] = 8'd120;
    sbox_22[194] = 8'd37;
    sbox_22[195] = 8'd46;
    sbox_22[196] = 8'd28;
    sbox_22[197] = 8'd166;
    sbox_22[198] = 8'd180;
    sbox_22[199] = 8'd198;
    sbox_22[200] = 8'd232;
    sbox_22[201] = 8'd221;
    sbox_22[202] = 8'd116;
    sbox_22[203] = 8'd31;
    sbox_22[204] = 8'd75;
    sbox_22[205] = 8'd189;
    sbox_22[206] = 8'd139;
    sbox_22[207] = 8'd138;
    sbox_22[208] = 8'd112;
    sbox_22[209] = 8'd62;
    sbox_22[210] = 8'd181;
    sbox_22[211] = 8'd102;
    sbox_22[212] = 8'd72;
    sbox_22[213] = 8'd3;
    sbox_22[214] = 8'd246;
    sbox_22[215] = 8'd14;
    sbox_22[216] = 8'd97;
    sbox_22[217] = 8'd53;
    sbox_22[218] = 8'd87;
    sbox_22[219] = 8'd185;
    sbox_22[220] = 8'd134;
    sbox_22[221] = 8'd193;
    sbox_22[222] = 8'd29;
    sbox_22[223] = 8'd158;
    sbox_22[224] = 8'd225;
    sbox_22[225] = 8'd248;
    sbox_22[226] = 8'd152;
    sbox_22[227] = 8'd17;
    sbox_22[228] = 8'd105;
    sbox_22[229] = 8'd217;
    sbox_22[230] = 8'd142;
    sbox_22[231] = 8'd148;
    sbox_22[232] = 8'd155;
    sbox_22[233] = 8'd30;
    sbox_22[234] = 8'd135;
    sbox_22[235] = 8'd233;
    sbox_22[236] = 8'd206;
    sbox_22[237] = 8'd85;
    sbox_22[238] = 8'd40;
    sbox_22[239] = 8'd223;
    sbox_22[240] = 8'd140;
    sbox_22[241] = 8'd161;
    sbox_22[242] = 8'd137;
    sbox_22[243] = 8'd13;
    sbox_22[244] = 8'd191;
    sbox_22[245] = 8'd230;
    sbox_22[246] = 8'd66;
    sbox_22[247] = 8'd104;
    sbox_22[248] = 8'd65;
    sbox_22[249] = 8'd153;
    sbox_22[250] = 8'd45;
    sbox_22[251] = 8'd15;
    sbox_22[252] = 8'd176;
    sbox_22[253] = 8'd84;
    sbox_22[254] = 8'd187;
    sbox_22[255] = 8'd22;
    sbox_23[0] = 8'd99;
    sbox_23[1] = 8'd124;
    sbox_23[2] = 8'd119;
    sbox_23[3] = 8'd123;
    sbox_23[4] = 8'd242;
    sbox_23[5] = 8'd107;
    sbox_23[6] = 8'd111;
    sbox_23[7] = 8'd197;
    sbox_23[8] = 8'd48;
    sbox_23[9] = 8'd1;
    sbox_23[10] = 8'd103;
    sbox_23[11] = 8'd43;
    sbox_23[12] = 8'd254;
    sbox_23[13] = 8'd215;
    sbox_23[14] = 8'd171;
    sbox_23[15] = 8'd118;
    sbox_23[16] = 8'd202;
    sbox_23[17] = 8'd130;
    sbox_23[18] = 8'd201;
    sbox_23[19] = 8'd125;
    sbox_23[20] = 8'd250;
    sbox_23[21] = 8'd89;
    sbox_23[22] = 8'd71;
    sbox_23[23] = 8'd240;
    sbox_23[24] = 8'd173;
    sbox_23[25] = 8'd212;
    sbox_23[26] = 8'd162;
    sbox_23[27] = 8'd175;
    sbox_23[28] = 8'd156;
    sbox_23[29] = 8'd164;
    sbox_23[30] = 8'd114;
    sbox_23[31] = 8'd192;
    sbox_23[32] = 8'd183;
    sbox_23[33] = 8'd253;
    sbox_23[34] = 8'd147;
    sbox_23[35] = 8'd38;
    sbox_23[36] = 8'd54;
    sbox_23[37] = 8'd63;
    sbox_23[38] = 8'd247;
    sbox_23[39] = 8'd204;
    sbox_23[40] = 8'd52;
    sbox_23[41] = 8'd165;
    sbox_23[42] = 8'd229;
    sbox_23[43] = 8'd241;
    sbox_23[44] = 8'd113;
    sbox_23[45] = 8'd216;
    sbox_23[46] = 8'd49;
    sbox_23[47] = 8'd21;
    sbox_23[48] = 8'd4;
    sbox_23[49] = 8'd199;
    sbox_23[50] = 8'd35;
    sbox_23[51] = 8'd195;
    sbox_23[52] = 8'd24;
    sbox_23[53] = 8'd150;
    sbox_23[54] = 8'd5;
    sbox_23[55] = 8'd154;
    sbox_23[56] = 8'd7;
    sbox_23[57] = 8'd18;
    sbox_23[58] = 8'd128;
    sbox_23[59] = 8'd226;
    sbox_23[60] = 8'd235;
    sbox_23[61] = 8'd39;
    sbox_23[62] = 8'd178;
    sbox_23[63] = 8'd117;
    sbox_23[64] = 8'd9;
    sbox_23[65] = 8'd131;
    sbox_23[66] = 8'd44;
    sbox_23[67] = 8'd26;
    sbox_23[68] = 8'd27;
    sbox_23[69] = 8'd110;
    sbox_23[70] = 8'd90;
    sbox_23[71] = 8'd160;
    sbox_23[72] = 8'd82;
    sbox_23[73] = 8'd59;
    sbox_23[74] = 8'd214;
    sbox_23[75] = 8'd179;
    sbox_23[76] = 8'd41;
    sbox_23[77] = 8'd227;
    sbox_23[78] = 8'd47;
    sbox_23[79] = 8'd132;
    sbox_23[80] = 8'd83;
    sbox_23[81] = 8'd209;
    sbox_23[82] = 8'd0;
    sbox_23[83] = 8'd237;
    sbox_23[84] = 8'd32;
    sbox_23[85] = 8'd252;
    sbox_23[86] = 8'd177;
    sbox_23[87] = 8'd91;
    sbox_23[88] = 8'd106;
    sbox_23[89] = 8'd203;
    sbox_23[90] = 8'd190;
    sbox_23[91] = 8'd57;
    sbox_23[92] = 8'd74;
    sbox_23[93] = 8'd76;
    sbox_23[94] = 8'd88;
    sbox_23[95] = 8'd207;
    sbox_23[96] = 8'd208;
    sbox_23[97] = 8'd239;
    sbox_23[98] = 8'd170;
    sbox_23[99] = 8'd251;
    sbox_23[100] = 8'd67;
    sbox_23[101] = 8'd77;
    sbox_23[102] = 8'd51;
    sbox_23[103] = 8'd133;
    sbox_23[104] = 8'd69;
    sbox_23[105] = 8'd249;
    sbox_23[106] = 8'd2;
    sbox_23[107] = 8'd127;
    sbox_23[108] = 8'd80;
    sbox_23[109] = 8'd60;
    sbox_23[110] = 8'd159;
    sbox_23[111] = 8'd168;
    sbox_23[112] = 8'd81;
    sbox_23[113] = 8'd163;
    sbox_23[114] = 8'd64;
    sbox_23[115] = 8'd143;
    sbox_23[116] = 8'd146;
    sbox_23[117] = 8'd157;
    sbox_23[118] = 8'd56;
    sbox_23[119] = 8'd245;
    sbox_23[120] = 8'd188;
    sbox_23[121] = 8'd182;
    sbox_23[122] = 8'd218;
    sbox_23[123] = 8'd33;
    sbox_23[124] = 8'd16;
    sbox_23[125] = 8'd255;
    sbox_23[126] = 8'd243;
    sbox_23[127] = 8'd210;
    sbox_23[128] = 8'd205;
    sbox_23[129] = 8'd12;
    sbox_23[130] = 8'd19;
    sbox_23[131] = 8'd236;
    sbox_23[132] = 8'd95;
    sbox_23[133] = 8'd151;
    sbox_23[134] = 8'd68;
    sbox_23[135] = 8'd23;
    sbox_23[136] = 8'd196;
    sbox_23[137] = 8'd167;
    sbox_23[138] = 8'd126;
    sbox_23[139] = 8'd61;
    sbox_23[140] = 8'd100;
    sbox_23[141] = 8'd93;
    sbox_23[142] = 8'd25;
    sbox_23[143] = 8'd115;
    sbox_23[144] = 8'd96;
    sbox_23[145] = 8'd129;
    sbox_23[146] = 8'd79;
    sbox_23[147] = 8'd220;
    sbox_23[148] = 8'd34;
    sbox_23[149] = 8'd42;
    sbox_23[150] = 8'd144;
    sbox_23[151] = 8'd136;
    sbox_23[152] = 8'd70;
    sbox_23[153] = 8'd238;
    sbox_23[154] = 8'd184;
    sbox_23[155] = 8'd20;
    sbox_23[156] = 8'd222;
    sbox_23[157] = 8'd94;
    sbox_23[158] = 8'd11;
    sbox_23[159] = 8'd219;
    sbox_23[160] = 8'd224;
    sbox_23[161] = 8'd50;
    sbox_23[162] = 8'd58;
    sbox_23[163] = 8'd10;
    sbox_23[164] = 8'd73;
    sbox_23[165] = 8'd6;
    sbox_23[166] = 8'd36;
    sbox_23[167] = 8'd92;
    sbox_23[168] = 8'd194;
    sbox_23[169] = 8'd211;
    sbox_23[170] = 8'd172;
    sbox_23[171] = 8'd98;
    sbox_23[172] = 8'd145;
    sbox_23[173] = 8'd149;
    sbox_23[174] = 8'd228;
    sbox_23[175] = 8'd121;
    sbox_23[176] = 8'd231;
    sbox_23[177] = 8'd200;
    sbox_23[178] = 8'd55;
    sbox_23[179] = 8'd109;
    sbox_23[180] = 8'd141;
    sbox_23[181] = 8'd213;
    sbox_23[182] = 8'd78;
    sbox_23[183] = 8'd169;
    sbox_23[184] = 8'd108;
    sbox_23[185] = 8'd86;
    sbox_23[186] = 8'd244;
    sbox_23[187] = 8'd234;
    sbox_23[188] = 8'd101;
    sbox_23[189] = 8'd122;
    sbox_23[190] = 8'd174;
    sbox_23[191] = 8'd8;
    sbox_23[192] = 8'd186;
    sbox_23[193] = 8'd120;
    sbox_23[194] = 8'd37;
    sbox_23[195] = 8'd46;
    sbox_23[196] = 8'd28;
    sbox_23[197] = 8'd166;
    sbox_23[198] = 8'd180;
    sbox_23[199] = 8'd198;
    sbox_23[200] = 8'd232;
    sbox_23[201] = 8'd221;
    sbox_23[202] = 8'd116;
    sbox_23[203] = 8'd31;
    sbox_23[204] = 8'd75;
    sbox_23[205] = 8'd189;
    sbox_23[206] = 8'd139;
    sbox_23[207] = 8'd138;
    sbox_23[208] = 8'd112;
    sbox_23[209] = 8'd62;
    sbox_23[210] = 8'd181;
    sbox_23[211] = 8'd102;
    sbox_23[212] = 8'd72;
    sbox_23[213] = 8'd3;
    sbox_23[214] = 8'd246;
    sbox_23[215] = 8'd14;
    sbox_23[216] = 8'd97;
    sbox_23[217] = 8'd53;
    sbox_23[218] = 8'd87;
    sbox_23[219] = 8'd185;
    sbox_23[220] = 8'd134;
    sbox_23[221] = 8'd193;
    sbox_23[222] = 8'd29;
    sbox_23[223] = 8'd158;
    sbox_23[224] = 8'd225;
    sbox_23[225] = 8'd248;
    sbox_23[226] = 8'd152;
    sbox_23[227] = 8'd17;
    sbox_23[228] = 8'd105;
    sbox_23[229] = 8'd217;
    sbox_23[230] = 8'd142;
    sbox_23[231] = 8'd148;
    sbox_23[232] = 8'd155;
    sbox_23[233] = 8'd30;
    sbox_23[234] = 8'd135;
    sbox_23[235] = 8'd233;
    sbox_23[236] = 8'd206;
    sbox_23[237] = 8'd85;
    sbox_23[238] = 8'd40;
    sbox_23[239] = 8'd223;
    sbox_23[240] = 8'd140;
    sbox_23[241] = 8'd161;
    sbox_23[242] = 8'd137;
    sbox_23[243] = 8'd13;
    sbox_23[244] = 8'd191;
    sbox_23[245] = 8'd230;
    sbox_23[246] = 8'd66;
    sbox_23[247] = 8'd104;
    sbox_23[248] = 8'd65;
    sbox_23[249] = 8'd153;
    sbox_23[250] = 8'd45;
    sbox_23[251] = 8'd15;
    sbox_23[252] = 8'd176;
    sbox_23[253] = 8'd84;
    sbox_23[254] = 8'd187;
    sbox_23[255] = 8'd22;
    sbox_24[0] = 8'd99;
    sbox_24[1] = 8'd124;
    sbox_24[2] = 8'd119;
    sbox_24[3] = 8'd123;
    sbox_24[4] = 8'd242;
    sbox_24[5] = 8'd107;
    sbox_24[6] = 8'd111;
    sbox_24[7] = 8'd197;
    sbox_24[8] = 8'd48;
    sbox_24[9] = 8'd1;
    sbox_24[10] = 8'd103;
    sbox_24[11] = 8'd43;
    sbox_24[12] = 8'd254;
    sbox_24[13] = 8'd215;
    sbox_24[14] = 8'd171;
    sbox_24[15] = 8'd118;
    sbox_24[16] = 8'd202;
    sbox_24[17] = 8'd130;
    sbox_24[18] = 8'd201;
    sbox_24[19] = 8'd125;
    sbox_24[20] = 8'd250;
    sbox_24[21] = 8'd89;
    sbox_24[22] = 8'd71;
    sbox_24[23] = 8'd240;
    sbox_24[24] = 8'd173;
    sbox_24[25] = 8'd212;
    sbox_24[26] = 8'd162;
    sbox_24[27] = 8'd175;
    sbox_24[28] = 8'd156;
    sbox_24[29] = 8'd164;
    sbox_24[30] = 8'd114;
    sbox_24[31] = 8'd192;
    sbox_24[32] = 8'd183;
    sbox_24[33] = 8'd253;
    sbox_24[34] = 8'd147;
    sbox_24[35] = 8'd38;
    sbox_24[36] = 8'd54;
    sbox_24[37] = 8'd63;
    sbox_24[38] = 8'd247;
    sbox_24[39] = 8'd204;
    sbox_24[40] = 8'd52;
    sbox_24[41] = 8'd165;
    sbox_24[42] = 8'd229;
    sbox_24[43] = 8'd241;
    sbox_24[44] = 8'd113;
    sbox_24[45] = 8'd216;
    sbox_24[46] = 8'd49;
    sbox_24[47] = 8'd21;
    sbox_24[48] = 8'd4;
    sbox_24[49] = 8'd199;
    sbox_24[50] = 8'd35;
    sbox_24[51] = 8'd195;
    sbox_24[52] = 8'd24;
    sbox_24[53] = 8'd150;
    sbox_24[54] = 8'd5;
    sbox_24[55] = 8'd154;
    sbox_24[56] = 8'd7;
    sbox_24[57] = 8'd18;
    sbox_24[58] = 8'd128;
    sbox_24[59] = 8'd226;
    sbox_24[60] = 8'd235;
    sbox_24[61] = 8'd39;
    sbox_24[62] = 8'd178;
    sbox_24[63] = 8'd117;
    sbox_24[64] = 8'd9;
    sbox_24[65] = 8'd131;
    sbox_24[66] = 8'd44;
    sbox_24[67] = 8'd26;
    sbox_24[68] = 8'd27;
    sbox_24[69] = 8'd110;
    sbox_24[70] = 8'd90;
    sbox_24[71] = 8'd160;
    sbox_24[72] = 8'd82;
    sbox_24[73] = 8'd59;
    sbox_24[74] = 8'd214;
    sbox_24[75] = 8'd179;
    sbox_24[76] = 8'd41;
    sbox_24[77] = 8'd227;
    sbox_24[78] = 8'd47;
    sbox_24[79] = 8'd132;
    sbox_24[80] = 8'd83;
    sbox_24[81] = 8'd209;
    sbox_24[82] = 8'd0;
    sbox_24[83] = 8'd237;
    sbox_24[84] = 8'd32;
    sbox_24[85] = 8'd252;
    sbox_24[86] = 8'd177;
    sbox_24[87] = 8'd91;
    sbox_24[88] = 8'd106;
    sbox_24[89] = 8'd203;
    sbox_24[90] = 8'd190;
    sbox_24[91] = 8'd57;
    sbox_24[92] = 8'd74;
    sbox_24[93] = 8'd76;
    sbox_24[94] = 8'd88;
    sbox_24[95] = 8'd207;
    sbox_24[96] = 8'd208;
    sbox_24[97] = 8'd239;
    sbox_24[98] = 8'd170;
    sbox_24[99] = 8'd251;
    sbox_24[100] = 8'd67;
    sbox_24[101] = 8'd77;
    sbox_24[102] = 8'd51;
    sbox_24[103] = 8'd133;
    sbox_24[104] = 8'd69;
    sbox_24[105] = 8'd249;
    sbox_24[106] = 8'd2;
    sbox_24[107] = 8'd127;
    sbox_24[108] = 8'd80;
    sbox_24[109] = 8'd60;
    sbox_24[110] = 8'd159;
    sbox_24[111] = 8'd168;
    sbox_24[112] = 8'd81;
    sbox_24[113] = 8'd163;
    sbox_24[114] = 8'd64;
    sbox_24[115] = 8'd143;
    sbox_24[116] = 8'd146;
    sbox_24[117] = 8'd157;
    sbox_24[118] = 8'd56;
    sbox_24[119] = 8'd245;
    sbox_24[120] = 8'd188;
    sbox_24[121] = 8'd182;
    sbox_24[122] = 8'd218;
    sbox_24[123] = 8'd33;
    sbox_24[124] = 8'd16;
    sbox_24[125] = 8'd255;
    sbox_24[126] = 8'd243;
    sbox_24[127] = 8'd210;
    sbox_24[128] = 8'd205;
    sbox_24[129] = 8'd12;
    sbox_24[130] = 8'd19;
    sbox_24[131] = 8'd236;
    sbox_24[132] = 8'd95;
    sbox_24[133] = 8'd151;
    sbox_24[134] = 8'd68;
    sbox_24[135] = 8'd23;
    sbox_24[136] = 8'd196;
    sbox_24[137] = 8'd167;
    sbox_24[138] = 8'd126;
    sbox_24[139] = 8'd61;
    sbox_24[140] = 8'd100;
    sbox_24[141] = 8'd93;
    sbox_24[142] = 8'd25;
    sbox_24[143] = 8'd115;
    sbox_24[144] = 8'd96;
    sbox_24[145] = 8'd129;
    sbox_24[146] = 8'd79;
    sbox_24[147] = 8'd220;
    sbox_24[148] = 8'd34;
    sbox_24[149] = 8'd42;
    sbox_24[150] = 8'd144;
    sbox_24[151] = 8'd136;
    sbox_24[152] = 8'd70;
    sbox_24[153] = 8'd238;
    sbox_24[154] = 8'd184;
    sbox_24[155] = 8'd20;
    sbox_24[156] = 8'd222;
    sbox_24[157] = 8'd94;
    sbox_24[158] = 8'd11;
    sbox_24[159] = 8'd219;
    sbox_24[160] = 8'd224;
    sbox_24[161] = 8'd50;
    sbox_24[162] = 8'd58;
    sbox_24[163] = 8'd10;
    sbox_24[164] = 8'd73;
    sbox_24[165] = 8'd6;
    sbox_24[166] = 8'd36;
    sbox_24[167] = 8'd92;
    sbox_24[168] = 8'd194;
    sbox_24[169] = 8'd211;
    sbox_24[170] = 8'd172;
    sbox_24[171] = 8'd98;
    sbox_24[172] = 8'd145;
    sbox_24[173] = 8'd149;
    sbox_24[174] = 8'd228;
    sbox_24[175] = 8'd121;
    sbox_24[176] = 8'd231;
    sbox_24[177] = 8'd200;
    sbox_24[178] = 8'd55;
    sbox_24[179] = 8'd109;
    sbox_24[180] = 8'd141;
    sbox_24[181] = 8'd213;
    sbox_24[182] = 8'd78;
    sbox_24[183] = 8'd169;
    sbox_24[184] = 8'd108;
    sbox_24[185] = 8'd86;
    sbox_24[186] = 8'd244;
    sbox_24[187] = 8'd234;
    sbox_24[188] = 8'd101;
    sbox_24[189] = 8'd122;
    sbox_24[190] = 8'd174;
    sbox_24[191] = 8'd8;
    sbox_24[192] = 8'd186;
    sbox_24[193] = 8'd120;
    sbox_24[194] = 8'd37;
    sbox_24[195] = 8'd46;
    sbox_24[196] = 8'd28;
    sbox_24[197] = 8'd166;
    sbox_24[198] = 8'd180;
    sbox_24[199] = 8'd198;
    sbox_24[200] = 8'd232;
    sbox_24[201] = 8'd221;
    sbox_24[202] = 8'd116;
    sbox_24[203] = 8'd31;
    sbox_24[204] = 8'd75;
    sbox_24[205] = 8'd189;
    sbox_24[206] = 8'd139;
    sbox_24[207] = 8'd138;
    sbox_24[208] = 8'd112;
    sbox_24[209] = 8'd62;
    sbox_24[210] = 8'd181;
    sbox_24[211] = 8'd102;
    sbox_24[212] = 8'd72;
    sbox_24[213] = 8'd3;
    sbox_24[214] = 8'd246;
    sbox_24[215] = 8'd14;
    sbox_24[216] = 8'd97;
    sbox_24[217] = 8'd53;
    sbox_24[218] = 8'd87;
    sbox_24[219] = 8'd185;
    sbox_24[220] = 8'd134;
    sbox_24[221] = 8'd193;
    sbox_24[222] = 8'd29;
    sbox_24[223] = 8'd158;
    sbox_24[224] = 8'd225;
    sbox_24[225] = 8'd248;
    sbox_24[226] = 8'd152;
    sbox_24[227] = 8'd17;
    sbox_24[228] = 8'd105;
    sbox_24[229] = 8'd217;
    sbox_24[230] = 8'd142;
    sbox_24[231] = 8'd148;
    sbox_24[232] = 8'd155;
    sbox_24[233] = 8'd30;
    sbox_24[234] = 8'd135;
    sbox_24[235] = 8'd233;
    sbox_24[236] = 8'd206;
    sbox_24[237] = 8'd85;
    sbox_24[238] = 8'd40;
    sbox_24[239] = 8'd223;
    sbox_24[240] = 8'd140;
    sbox_24[241] = 8'd161;
    sbox_24[242] = 8'd137;
    sbox_24[243] = 8'd13;
    sbox_24[244] = 8'd191;
    sbox_24[245] = 8'd230;
    sbox_24[246] = 8'd66;
    sbox_24[247] = 8'd104;
    sbox_24[248] = 8'd65;
    sbox_24[249] = 8'd153;
    sbox_24[250] = 8'd45;
    sbox_24[251] = 8'd15;
    sbox_24[252] = 8'd176;
    sbox_24[253] = 8'd84;
    sbox_24[254] = 8'd187;
    sbox_24[255] = 8'd22;
    sbox_25[0] = 8'd99;
    sbox_25[1] = 8'd124;
    sbox_25[2] = 8'd119;
    sbox_25[3] = 8'd123;
    sbox_25[4] = 8'd242;
    sbox_25[5] = 8'd107;
    sbox_25[6] = 8'd111;
    sbox_25[7] = 8'd197;
    sbox_25[8] = 8'd48;
    sbox_25[9] = 8'd1;
    sbox_25[10] = 8'd103;
    sbox_25[11] = 8'd43;
    sbox_25[12] = 8'd254;
    sbox_25[13] = 8'd215;
    sbox_25[14] = 8'd171;
    sbox_25[15] = 8'd118;
    sbox_25[16] = 8'd202;
    sbox_25[17] = 8'd130;
    sbox_25[18] = 8'd201;
    sbox_25[19] = 8'd125;
    sbox_25[20] = 8'd250;
    sbox_25[21] = 8'd89;
    sbox_25[22] = 8'd71;
    sbox_25[23] = 8'd240;
    sbox_25[24] = 8'd173;
    sbox_25[25] = 8'd212;
    sbox_25[26] = 8'd162;
    sbox_25[27] = 8'd175;
    sbox_25[28] = 8'd156;
    sbox_25[29] = 8'd164;
    sbox_25[30] = 8'd114;
    sbox_25[31] = 8'd192;
    sbox_25[32] = 8'd183;
    sbox_25[33] = 8'd253;
    sbox_25[34] = 8'd147;
    sbox_25[35] = 8'd38;
    sbox_25[36] = 8'd54;
    sbox_25[37] = 8'd63;
    sbox_25[38] = 8'd247;
    sbox_25[39] = 8'd204;
    sbox_25[40] = 8'd52;
    sbox_25[41] = 8'd165;
    sbox_25[42] = 8'd229;
    sbox_25[43] = 8'd241;
    sbox_25[44] = 8'd113;
    sbox_25[45] = 8'd216;
    sbox_25[46] = 8'd49;
    sbox_25[47] = 8'd21;
    sbox_25[48] = 8'd4;
    sbox_25[49] = 8'd199;
    sbox_25[50] = 8'd35;
    sbox_25[51] = 8'd195;
    sbox_25[52] = 8'd24;
    sbox_25[53] = 8'd150;
    sbox_25[54] = 8'd5;
    sbox_25[55] = 8'd154;
    sbox_25[56] = 8'd7;
    sbox_25[57] = 8'd18;
    sbox_25[58] = 8'd128;
    sbox_25[59] = 8'd226;
    sbox_25[60] = 8'd235;
    sbox_25[61] = 8'd39;
    sbox_25[62] = 8'd178;
    sbox_25[63] = 8'd117;
    sbox_25[64] = 8'd9;
    sbox_25[65] = 8'd131;
    sbox_25[66] = 8'd44;
    sbox_25[67] = 8'd26;
    sbox_25[68] = 8'd27;
    sbox_25[69] = 8'd110;
    sbox_25[70] = 8'd90;
    sbox_25[71] = 8'd160;
    sbox_25[72] = 8'd82;
    sbox_25[73] = 8'd59;
    sbox_25[74] = 8'd214;
    sbox_25[75] = 8'd179;
    sbox_25[76] = 8'd41;
    sbox_25[77] = 8'd227;
    sbox_25[78] = 8'd47;
    sbox_25[79] = 8'd132;
    sbox_25[80] = 8'd83;
    sbox_25[81] = 8'd209;
    sbox_25[82] = 8'd0;
    sbox_25[83] = 8'd237;
    sbox_25[84] = 8'd32;
    sbox_25[85] = 8'd252;
    sbox_25[86] = 8'd177;
    sbox_25[87] = 8'd91;
    sbox_25[88] = 8'd106;
    sbox_25[89] = 8'd203;
    sbox_25[90] = 8'd190;
    sbox_25[91] = 8'd57;
    sbox_25[92] = 8'd74;
    sbox_25[93] = 8'd76;
    sbox_25[94] = 8'd88;
    sbox_25[95] = 8'd207;
    sbox_25[96] = 8'd208;
    sbox_25[97] = 8'd239;
    sbox_25[98] = 8'd170;
    sbox_25[99] = 8'd251;
    sbox_25[100] = 8'd67;
    sbox_25[101] = 8'd77;
    sbox_25[102] = 8'd51;
    sbox_25[103] = 8'd133;
    sbox_25[104] = 8'd69;
    sbox_25[105] = 8'd249;
    sbox_25[106] = 8'd2;
    sbox_25[107] = 8'd127;
    sbox_25[108] = 8'd80;
    sbox_25[109] = 8'd60;
    sbox_25[110] = 8'd159;
    sbox_25[111] = 8'd168;
    sbox_25[112] = 8'd81;
    sbox_25[113] = 8'd163;
    sbox_25[114] = 8'd64;
    sbox_25[115] = 8'd143;
    sbox_25[116] = 8'd146;
    sbox_25[117] = 8'd157;
    sbox_25[118] = 8'd56;
    sbox_25[119] = 8'd245;
    sbox_25[120] = 8'd188;
    sbox_25[121] = 8'd182;
    sbox_25[122] = 8'd218;
    sbox_25[123] = 8'd33;
    sbox_25[124] = 8'd16;
    sbox_25[125] = 8'd255;
    sbox_25[126] = 8'd243;
    sbox_25[127] = 8'd210;
    sbox_25[128] = 8'd205;
    sbox_25[129] = 8'd12;
    sbox_25[130] = 8'd19;
    sbox_25[131] = 8'd236;
    sbox_25[132] = 8'd95;
    sbox_25[133] = 8'd151;
    sbox_25[134] = 8'd68;
    sbox_25[135] = 8'd23;
    sbox_25[136] = 8'd196;
    sbox_25[137] = 8'd167;
    sbox_25[138] = 8'd126;
    sbox_25[139] = 8'd61;
    sbox_25[140] = 8'd100;
    sbox_25[141] = 8'd93;
    sbox_25[142] = 8'd25;
    sbox_25[143] = 8'd115;
    sbox_25[144] = 8'd96;
    sbox_25[145] = 8'd129;
    sbox_25[146] = 8'd79;
    sbox_25[147] = 8'd220;
    sbox_25[148] = 8'd34;
    sbox_25[149] = 8'd42;
    sbox_25[150] = 8'd144;
    sbox_25[151] = 8'd136;
    sbox_25[152] = 8'd70;
    sbox_25[153] = 8'd238;
    sbox_25[154] = 8'd184;
    sbox_25[155] = 8'd20;
    sbox_25[156] = 8'd222;
    sbox_25[157] = 8'd94;
    sbox_25[158] = 8'd11;
    sbox_25[159] = 8'd219;
    sbox_25[160] = 8'd224;
    sbox_25[161] = 8'd50;
    sbox_25[162] = 8'd58;
    sbox_25[163] = 8'd10;
    sbox_25[164] = 8'd73;
    sbox_25[165] = 8'd6;
    sbox_25[166] = 8'd36;
    sbox_25[167] = 8'd92;
    sbox_25[168] = 8'd194;
    sbox_25[169] = 8'd211;
    sbox_25[170] = 8'd172;
    sbox_25[171] = 8'd98;
    sbox_25[172] = 8'd145;
    sbox_25[173] = 8'd149;
    sbox_25[174] = 8'd228;
    sbox_25[175] = 8'd121;
    sbox_25[176] = 8'd231;
    sbox_25[177] = 8'd200;
    sbox_25[178] = 8'd55;
    sbox_25[179] = 8'd109;
    sbox_25[180] = 8'd141;
    sbox_25[181] = 8'd213;
    sbox_25[182] = 8'd78;
    sbox_25[183] = 8'd169;
    sbox_25[184] = 8'd108;
    sbox_25[185] = 8'd86;
    sbox_25[186] = 8'd244;
    sbox_25[187] = 8'd234;
    sbox_25[188] = 8'd101;
    sbox_25[189] = 8'd122;
    sbox_25[190] = 8'd174;
    sbox_25[191] = 8'd8;
    sbox_25[192] = 8'd186;
    sbox_25[193] = 8'd120;
    sbox_25[194] = 8'd37;
    sbox_25[195] = 8'd46;
    sbox_25[196] = 8'd28;
    sbox_25[197] = 8'd166;
    sbox_25[198] = 8'd180;
    sbox_25[199] = 8'd198;
    sbox_25[200] = 8'd232;
    sbox_25[201] = 8'd221;
    sbox_25[202] = 8'd116;
    sbox_25[203] = 8'd31;
    sbox_25[204] = 8'd75;
    sbox_25[205] = 8'd189;
    sbox_25[206] = 8'd139;
    sbox_25[207] = 8'd138;
    sbox_25[208] = 8'd112;
    sbox_25[209] = 8'd62;
    sbox_25[210] = 8'd181;
    sbox_25[211] = 8'd102;
    sbox_25[212] = 8'd72;
    sbox_25[213] = 8'd3;
    sbox_25[214] = 8'd246;
    sbox_25[215] = 8'd14;
    sbox_25[216] = 8'd97;
    sbox_25[217] = 8'd53;
    sbox_25[218] = 8'd87;
    sbox_25[219] = 8'd185;
    sbox_25[220] = 8'd134;
    sbox_25[221] = 8'd193;
    sbox_25[222] = 8'd29;
    sbox_25[223] = 8'd158;
    sbox_25[224] = 8'd225;
    sbox_25[225] = 8'd248;
    sbox_25[226] = 8'd152;
    sbox_25[227] = 8'd17;
    sbox_25[228] = 8'd105;
    sbox_25[229] = 8'd217;
    sbox_25[230] = 8'd142;
    sbox_25[231] = 8'd148;
    sbox_25[232] = 8'd155;
    sbox_25[233] = 8'd30;
    sbox_25[234] = 8'd135;
    sbox_25[235] = 8'd233;
    sbox_25[236] = 8'd206;
    sbox_25[237] = 8'd85;
    sbox_25[238] = 8'd40;
    sbox_25[239] = 8'd223;
    sbox_25[240] = 8'd140;
    sbox_25[241] = 8'd161;
    sbox_25[242] = 8'd137;
    sbox_25[243] = 8'd13;
    sbox_25[244] = 8'd191;
    sbox_25[245] = 8'd230;
    sbox_25[246] = 8'd66;
    sbox_25[247] = 8'd104;
    sbox_25[248] = 8'd65;
    sbox_25[249] = 8'd153;
    sbox_25[250] = 8'd45;
    sbox_25[251] = 8'd15;
    sbox_25[252] = 8'd176;
    sbox_25[253] = 8'd84;
    sbox_25[254] = 8'd187;
    sbox_25[255] = 8'd22;
    sbox_26[0] = 8'd99;
    sbox_26[1] = 8'd124;
    sbox_26[2] = 8'd119;
    sbox_26[3] = 8'd123;
    sbox_26[4] = 8'd242;
    sbox_26[5] = 8'd107;
    sbox_26[6] = 8'd111;
    sbox_26[7] = 8'd197;
    sbox_26[8] = 8'd48;
    sbox_26[9] = 8'd1;
    sbox_26[10] = 8'd103;
    sbox_26[11] = 8'd43;
    sbox_26[12] = 8'd254;
    sbox_26[13] = 8'd215;
    sbox_26[14] = 8'd171;
    sbox_26[15] = 8'd118;
    sbox_26[16] = 8'd202;
    sbox_26[17] = 8'd130;
    sbox_26[18] = 8'd201;
    sbox_26[19] = 8'd125;
    sbox_26[20] = 8'd250;
    sbox_26[21] = 8'd89;
    sbox_26[22] = 8'd71;
    sbox_26[23] = 8'd240;
    sbox_26[24] = 8'd173;
    sbox_26[25] = 8'd212;
    sbox_26[26] = 8'd162;
    sbox_26[27] = 8'd175;
    sbox_26[28] = 8'd156;
    sbox_26[29] = 8'd164;
    sbox_26[30] = 8'd114;
    sbox_26[31] = 8'd192;
    sbox_26[32] = 8'd183;
    sbox_26[33] = 8'd253;
    sbox_26[34] = 8'd147;
    sbox_26[35] = 8'd38;
    sbox_26[36] = 8'd54;
    sbox_26[37] = 8'd63;
    sbox_26[38] = 8'd247;
    sbox_26[39] = 8'd204;
    sbox_26[40] = 8'd52;
    sbox_26[41] = 8'd165;
    sbox_26[42] = 8'd229;
    sbox_26[43] = 8'd241;
    sbox_26[44] = 8'd113;
    sbox_26[45] = 8'd216;
    sbox_26[46] = 8'd49;
    sbox_26[47] = 8'd21;
    sbox_26[48] = 8'd4;
    sbox_26[49] = 8'd199;
    sbox_26[50] = 8'd35;
    sbox_26[51] = 8'd195;
    sbox_26[52] = 8'd24;
    sbox_26[53] = 8'd150;
    sbox_26[54] = 8'd5;
    sbox_26[55] = 8'd154;
    sbox_26[56] = 8'd7;
    sbox_26[57] = 8'd18;
    sbox_26[58] = 8'd128;
    sbox_26[59] = 8'd226;
    sbox_26[60] = 8'd235;
    sbox_26[61] = 8'd39;
    sbox_26[62] = 8'd178;
    sbox_26[63] = 8'd117;
    sbox_26[64] = 8'd9;
    sbox_26[65] = 8'd131;
    sbox_26[66] = 8'd44;
    sbox_26[67] = 8'd26;
    sbox_26[68] = 8'd27;
    sbox_26[69] = 8'd110;
    sbox_26[70] = 8'd90;
    sbox_26[71] = 8'd160;
    sbox_26[72] = 8'd82;
    sbox_26[73] = 8'd59;
    sbox_26[74] = 8'd214;
    sbox_26[75] = 8'd179;
    sbox_26[76] = 8'd41;
    sbox_26[77] = 8'd227;
    sbox_26[78] = 8'd47;
    sbox_26[79] = 8'd132;
    sbox_26[80] = 8'd83;
    sbox_26[81] = 8'd209;
    sbox_26[82] = 8'd0;
    sbox_26[83] = 8'd237;
    sbox_26[84] = 8'd32;
    sbox_26[85] = 8'd252;
    sbox_26[86] = 8'd177;
    sbox_26[87] = 8'd91;
    sbox_26[88] = 8'd106;
    sbox_26[89] = 8'd203;
    sbox_26[90] = 8'd190;
    sbox_26[91] = 8'd57;
    sbox_26[92] = 8'd74;
    sbox_26[93] = 8'd76;
    sbox_26[94] = 8'd88;
    sbox_26[95] = 8'd207;
    sbox_26[96] = 8'd208;
    sbox_26[97] = 8'd239;
    sbox_26[98] = 8'd170;
    sbox_26[99] = 8'd251;
    sbox_26[100] = 8'd67;
    sbox_26[101] = 8'd77;
    sbox_26[102] = 8'd51;
    sbox_26[103] = 8'd133;
    sbox_26[104] = 8'd69;
    sbox_26[105] = 8'd249;
    sbox_26[106] = 8'd2;
    sbox_26[107] = 8'd127;
    sbox_26[108] = 8'd80;
    sbox_26[109] = 8'd60;
    sbox_26[110] = 8'd159;
    sbox_26[111] = 8'd168;
    sbox_26[112] = 8'd81;
    sbox_26[113] = 8'd163;
    sbox_26[114] = 8'd64;
    sbox_26[115] = 8'd143;
    sbox_26[116] = 8'd146;
    sbox_26[117] = 8'd157;
    sbox_26[118] = 8'd56;
    sbox_26[119] = 8'd245;
    sbox_26[120] = 8'd188;
    sbox_26[121] = 8'd182;
    sbox_26[122] = 8'd218;
    sbox_26[123] = 8'd33;
    sbox_26[124] = 8'd16;
    sbox_26[125] = 8'd255;
    sbox_26[126] = 8'd243;
    sbox_26[127] = 8'd210;
    sbox_26[128] = 8'd205;
    sbox_26[129] = 8'd12;
    sbox_26[130] = 8'd19;
    sbox_26[131] = 8'd236;
    sbox_26[132] = 8'd95;
    sbox_26[133] = 8'd151;
    sbox_26[134] = 8'd68;
    sbox_26[135] = 8'd23;
    sbox_26[136] = 8'd196;
    sbox_26[137] = 8'd167;
    sbox_26[138] = 8'd126;
    sbox_26[139] = 8'd61;
    sbox_26[140] = 8'd100;
    sbox_26[141] = 8'd93;
    sbox_26[142] = 8'd25;
    sbox_26[143] = 8'd115;
    sbox_26[144] = 8'd96;
    sbox_26[145] = 8'd129;
    sbox_26[146] = 8'd79;
    sbox_26[147] = 8'd220;
    sbox_26[148] = 8'd34;
    sbox_26[149] = 8'd42;
    sbox_26[150] = 8'd144;
    sbox_26[151] = 8'd136;
    sbox_26[152] = 8'd70;
    sbox_26[153] = 8'd238;
    sbox_26[154] = 8'd184;
    sbox_26[155] = 8'd20;
    sbox_26[156] = 8'd222;
    sbox_26[157] = 8'd94;
    sbox_26[158] = 8'd11;
    sbox_26[159] = 8'd219;
    sbox_26[160] = 8'd224;
    sbox_26[161] = 8'd50;
    sbox_26[162] = 8'd58;
    sbox_26[163] = 8'd10;
    sbox_26[164] = 8'd73;
    sbox_26[165] = 8'd6;
    sbox_26[166] = 8'd36;
    sbox_26[167] = 8'd92;
    sbox_26[168] = 8'd194;
    sbox_26[169] = 8'd211;
    sbox_26[170] = 8'd172;
    sbox_26[171] = 8'd98;
    sbox_26[172] = 8'd145;
    sbox_26[173] = 8'd149;
    sbox_26[174] = 8'd228;
    sbox_26[175] = 8'd121;
    sbox_26[176] = 8'd231;
    sbox_26[177] = 8'd200;
    sbox_26[178] = 8'd55;
    sbox_26[179] = 8'd109;
    sbox_26[180] = 8'd141;
    sbox_26[181] = 8'd213;
    sbox_26[182] = 8'd78;
    sbox_26[183] = 8'd169;
    sbox_26[184] = 8'd108;
    sbox_26[185] = 8'd86;
    sbox_26[186] = 8'd244;
    sbox_26[187] = 8'd234;
    sbox_26[188] = 8'd101;
    sbox_26[189] = 8'd122;
    sbox_26[190] = 8'd174;
    sbox_26[191] = 8'd8;
    sbox_26[192] = 8'd186;
    sbox_26[193] = 8'd120;
    sbox_26[194] = 8'd37;
    sbox_26[195] = 8'd46;
    sbox_26[196] = 8'd28;
    sbox_26[197] = 8'd166;
    sbox_26[198] = 8'd180;
    sbox_26[199] = 8'd198;
    sbox_26[200] = 8'd232;
    sbox_26[201] = 8'd221;
    sbox_26[202] = 8'd116;
    sbox_26[203] = 8'd31;
    sbox_26[204] = 8'd75;
    sbox_26[205] = 8'd189;
    sbox_26[206] = 8'd139;
    sbox_26[207] = 8'd138;
    sbox_26[208] = 8'd112;
    sbox_26[209] = 8'd62;
    sbox_26[210] = 8'd181;
    sbox_26[211] = 8'd102;
    sbox_26[212] = 8'd72;
    sbox_26[213] = 8'd3;
    sbox_26[214] = 8'd246;
    sbox_26[215] = 8'd14;
    sbox_26[216] = 8'd97;
    sbox_26[217] = 8'd53;
    sbox_26[218] = 8'd87;
    sbox_26[219] = 8'd185;
    sbox_26[220] = 8'd134;
    sbox_26[221] = 8'd193;
    sbox_26[222] = 8'd29;
    sbox_26[223] = 8'd158;
    sbox_26[224] = 8'd225;
    sbox_26[225] = 8'd248;
    sbox_26[226] = 8'd152;
    sbox_26[227] = 8'd17;
    sbox_26[228] = 8'd105;
    sbox_26[229] = 8'd217;
    sbox_26[230] = 8'd142;
    sbox_26[231] = 8'd148;
    sbox_26[232] = 8'd155;
    sbox_26[233] = 8'd30;
    sbox_26[234] = 8'd135;
    sbox_26[235] = 8'd233;
    sbox_26[236] = 8'd206;
    sbox_26[237] = 8'd85;
    sbox_26[238] = 8'd40;
    sbox_26[239] = 8'd223;
    sbox_26[240] = 8'd140;
    sbox_26[241] = 8'd161;
    sbox_26[242] = 8'd137;
    sbox_26[243] = 8'd13;
    sbox_26[244] = 8'd191;
    sbox_26[245] = 8'd230;
    sbox_26[246] = 8'd66;
    sbox_26[247] = 8'd104;
    sbox_26[248] = 8'd65;
    sbox_26[249] = 8'd153;
    sbox_26[250] = 8'd45;
    sbox_26[251] = 8'd15;
    sbox_26[252] = 8'd176;
    sbox_26[253] = 8'd84;
    sbox_26[254] = 8'd187;
    sbox_26[255] = 8'd22;
    sbox_27[0] = 8'd99;
    sbox_27[1] = 8'd124;
    sbox_27[2] = 8'd119;
    sbox_27[3] = 8'd123;
    sbox_27[4] = 8'd242;
    sbox_27[5] = 8'd107;
    sbox_27[6] = 8'd111;
    sbox_27[7] = 8'd197;
    sbox_27[8] = 8'd48;
    sbox_27[9] = 8'd1;
    sbox_27[10] = 8'd103;
    sbox_27[11] = 8'd43;
    sbox_27[12] = 8'd254;
    sbox_27[13] = 8'd215;
    sbox_27[14] = 8'd171;
    sbox_27[15] = 8'd118;
    sbox_27[16] = 8'd202;
    sbox_27[17] = 8'd130;
    sbox_27[18] = 8'd201;
    sbox_27[19] = 8'd125;
    sbox_27[20] = 8'd250;
    sbox_27[21] = 8'd89;
    sbox_27[22] = 8'd71;
    sbox_27[23] = 8'd240;
    sbox_27[24] = 8'd173;
    sbox_27[25] = 8'd212;
    sbox_27[26] = 8'd162;
    sbox_27[27] = 8'd175;
    sbox_27[28] = 8'd156;
    sbox_27[29] = 8'd164;
    sbox_27[30] = 8'd114;
    sbox_27[31] = 8'd192;
    sbox_27[32] = 8'd183;
    sbox_27[33] = 8'd253;
    sbox_27[34] = 8'd147;
    sbox_27[35] = 8'd38;
    sbox_27[36] = 8'd54;
    sbox_27[37] = 8'd63;
    sbox_27[38] = 8'd247;
    sbox_27[39] = 8'd204;
    sbox_27[40] = 8'd52;
    sbox_27[41] = 8'd165;
    sbox_27[42] = 8'd229;
    sbox_27[43] = 8'd241;
    sbox_27[44] = 8'd113;
    sbox_27[45] = 8'd216;
    sbox_27[46] = 8'd49;
    sbox_27[47] = 8'd21;
    sbox_27[48] = 8'd4;
    sbox_27[49] = 8'd199;
    sbox_27[50] = 8'd35;
    sbox_27[51] = 8'd195;
    sbox_27[52] = 8'd24;
    sbox_27[53] = 8'd150;
    sbox_27[54] = 8'd5;
    sbox_27[55] = 8'd154;
    sbox_27[56] = 8'd7;
    sbox_27[57] = 8'd18;
    sbox_27[58] = 8'd128;
    sbox_27[59] = 8'd226;
    sbox_27[60] = 8'd235;
    sbox_27[61] = 8'd39;
    sbox_27[62] = 8'd178;
    sbox_27[63] = 8'd117;
    sbox_27[64] = 8'd9;
    sbox_27[65] = 8'd131;
    sbox_27[66] = 8'd44;
    sbox_27[67] = 8'd26;
    sbox_27[68] = 8'd27;
    sbox_27[69] = 8'd110;
    sbox_27[70] = 8'd90;
    sbox_27[71] = 8'd160;
    sbox_27[72] = 8'd82;
    sbox_27[73] = 8'd59;
    sbox_27[74] = 8'd214;
    sbox_27[75] = 8'd179;
    sbox_27[76] = 8'd41;
    sbox_27[77] = 8'd227;
    sbox_27[78] = 8'd47;
    sbox_27[79] = 8'd132;
    sbox_27[80] = 8'd83;
    sbox_27[81] = 8'd209;
    sbox_27[82] = 8'd0;
    sbox_27[83] = 8'd237;
    sbox_27[84] = 8'd32;
    sbox_27[85] = 8'd252;
    sbox_27[86] = 8'd177;
    sbox_27[87] = 8'd91;
    sbox_27[88] = 8'd106;
    sbox_27[89] = 8'd203;
    sbox_27[90] = 8'd190;
    sbox_27[91] = 8'd57;
    sbox_27[92] = 8'd74;
    sbox_27[93] = 8'd76;
    sbox_27[94] = 8'd88;
    sbox_27[95] = 8'd207;
    sbox_27[96] = 8'd208;
    sbox_27[97] = 8'd239;
    sbox_27[98] = 8'd170;
    sbox_27[99] = 8'd251;
    sbox_27[100] = 8'd67;
    sbox_27[101] = 8'd77;
    sbox_27[102] = 8'd51;
    sbox_27[103] = 8'd133;
    sbox_27[104] = 8'd69;
    sbox_27[105] = 8'd249;
    sbox_27[106] = 8'd2;
    sbox_27[107] = 8'd127;
    sbox_27[108] = 8'd80;
    sbox_27[109] = 8'd60;
    sbox_27[110] = 8'd159;
    sbox_27[111] = 8'd168;
    sbox_27[112] = 8'd81;
    sbox_27[113] = 8'd163;
    sbox_27[114] = 8'd64;
    sbox_27[115] = 8'd143;
    sbox_27[116] = 8'd146;
    sbox_27[117] = 8'd157;
    sbox_27[118] = 8'd56;
    sbox_27[119] = 8'd245;
    sbox_27[120] = 8'd188;
    sbox_27[121] = 8'd182;
    sbox_27[122] = 8'd218;
    sbox_27[123] = 8'd33;
    sbox_27[124] = 8'd16;
    sbox_27[125] = 8'd255;
    sbox_27[126] = 8'd243;
    sbox_27[127] = 8'd210;
    sbox_27[128] = 8'd205;
    sbox_27[129] = 8'd12;
    sbox_27[130] = 8'd19;
    sbox_27[131] = 8'd236;
    sbox_27[132] = 8'd95;
    sbox_27[133] = 8'd151;
    sbox_27[134] = 8'd68;
    sbox_27[135] = 8'd23;
    sbox_27[136] = 8'd196;
    sbox_27[137] = 8'd167;
    sbox_27[138] = 8'd126;
    sbox_27[139] = 8'd61;
    sbox_27[140] = 8'd100;
    sbox_27[141] = 8'd93;
    sbox_27[142] = 8'd25;
    sbox_27[143] = 8'd115;
    sbox_27[144] = 8'd96;
    sbox_27[145] = 8'd129;
    sbox_27[146] = 8'd79;
    sbox_27[147] = 8'd220;
    sbox_27[148] = 8'd34;
    sbox_27[149] = 8'd42;
    sbox_27[150] = 8'd144;
    sbox_27[151] = 8'd136;
    sbox_27[152] = 8'd70;
    sbox_27[153] = 8'd238;
    sbox_27[154] = 8'd184;
    sbox_27[155] = 8'd20;
    sbox_27[156] = 8'd222;
    sbox_27[157] = 8'd94;
    sbox_27[158] = 8'd11;
    sbox_27[159] = 8'd219;
    sbox_27[160] = 8'd224;
    sbox_27[161] = 8'd50;
    sbox_27[162] = 8'd58;
    sbox_27[163] = 8'd10;
    sbox_27[164] = 8'd73;
    sbox_27[165] = 8'd6;
    sbox_27[166] = 8'd36;
    sbox_27[167] = 8'd92;
    sbox_27[168] = 8'd194;
    sbox_27[169] = 8'd211;
    sbox_27[170] = 8'd172;
    sbox_27[171] = 8'd98;
    sbox_27[172] = 8'd145;
    sbox_27[173] = 8'd149;
    sbox_27[174] = 8'd228;
    sbox_27[175] = 8'd121;
    sbox_27[176] = 8'd231;
    sbox_27[177] = 8'd200;
    sbox_27[178] = 8'd55;
    sbox_27[179] = 8'd109;
    sbox_27[180] = 8'd141;
    sbox_27[181] = 8'd213;
    sbox_27[182] = 8'd78;
    sbox_27[183] = 8'd169;
    sbox_27[184] = 8'd108;
    sbox_27[185] = 8'd86;
    sbox_27[186] = 8'd244;
    sbox_27[187] = 8'd234;
    sbox_27[188] = 8'd101;
    sbox_27[189] = 8'd122;
    sbox_27[190] = 8'd174;
    sbox_27[191] = 8'd8;
    sbox_27[192] = 8'd186;
    sbox_27[193] = 8'd120;
    sbox_27[194] = 8'd37;
    sbox_27[195] = 8'd46;
    sbox_27[196] = 8'd28;
    sbox_27[197] = 8'd166;
    sbox_27[198] = 8'd180;
    sbox_27[199] = 8'd198;
    sbox_27[200] = 8'd232;
    sbox_27[201] = 8'd221;
    sbox_27[202] = 8'd116;
    sbox_27[203] = 8'd31;
    sbox_27[204] = 8'd75;
    sbox_27[205] = 8'd189;
    sbox_27[206] = 8'd139;
    sbox_27[207] = 8'd138;
    sbox_27[208] = 8'd112;
    sbox_27[209] = 8'd62;
    sbox_27[210] = 8'd181;
    sbox_27[211] = 8'd102;
    sbox_27[212] = 8'd72;
    sbox_27[213] = 8'd3;
    sbox_27[214] = 8'd246;
    sbox_27[215] = 8'd14;
    sbox_27[216] = 8'd97;
    sbox_27[217] = 8'd53;
    sbox_27[218] = 8'd87;
    sbox_27[219] = 8'd185;
    sbox_27[220] = 8'd134;
    sbox_27[221] = 8'd193;
    sbox_27[222] = 8'd29;
    sbox_27[223] = 8'd158;
    sbox_27[224] = 8'd225;
    sbox_27[225] = 8'd248;
    sbox_27[226] = 8'd152;
    sbox_27[227] = 8'd17;
    sbox_27[228] = 8'd105;
    sbox_27[229] = 8'd217;
    sbox_27[230] = 8'd142;
    sbox_27[231] = 8'd148;
    sbox_27[232] = 8'd155;
    sbox_27[233] = 8'd30;
    sbox_27[234] = 8'd135;
    sbox_27[235] = 8'd233;
    sbox_27[236] = 8'd206;
    sbox_27[237] = 8'd85;
    sbox_27[238] = 8'd40;
    sbox_27[239] = 8'd223;
    sbox_27[240] = 8'd140;
    sbox_27[241] = 8'd161;
    sbox_27[242] = 8'd137;
    sbox_27[243] = 8'd13;
    sbox_27[244] = 8'd191;
    sbox_27[245] = 8'd230;
    sbox_27[246] = 8'd66;
    sbox_27[247] = 8'd104;
    sbox_27[248] = 8'd65;
    sbox_27[249] = 8'd153;
    sbox_27[250] = 8'd45;
    sbox_27[251] = 8'd15;
    sbox_27[252] = 8'd176;
    sbox_27[253] = 8'd84;
    sbox_27[254] = 8'd187;
    sbox_27[255] = 8'd22;
    sbox_28[0] = 8'd99;
    sbox_28[1] = 8'd124;
    sbox_28[2] = 8'd119;
    sbox_28[3] = 8'd123;
    sbox_28[4] = 8'd242;
    sbox_28[5] = 8'd107;
    sbox_28[6] = 8'd111;
    sbox_28[7] = 8'd197;
    sbox_28[8] = 8'd48;
    sbox_28[9] = 8'd1;
    sbox_28[10] = 8'd103;
    sbox_28[11] = 8'd43;
    sbox_28[12] = 8'd254;
    sbox_28[13] = 8'd215;
    sbox_28[14] = 8'd171;
    sbox_28[15] = 8'd118;
    sbox_28[16] = 8'd202;
    sbox_28[17] = 8'd130;
    sbox_28[18] = 8'd201;
    sbox_28[19] = 8'd125;
    sbox_28[20] = 8'd250;
    sbox_28[21] = 8'd89;
    sbox_28[22] = 8'd71;
    sbox_28[23] = 8'd240;
    sbox_28[24] = 8'd173;
    sbox_28[25] = 8'd212;
    sbox_28[26] = 8'd162;
    sbox_28[27] = 8'd175;
    sbox_28[28] = 8'd156;
    sbox_28[29] = 8'd164;
    sbox_28[30] = 8'd114;
    sbox_28[31] = 8'd192;
    sbox_28[32] = 8'd183;
    sbox_28[33] = 8'd253;
    sbox_28[34] = 8'd147;
    sbox_28[35] = 8'd38;
    sbox_28[36] = 8'd54;
    sbox_28[37] = 8'd63;
    sbox_28[38] = 8'd247;
    sbox_28[39] = 8'd204;
    sbox_28[40] = 8'd52;
    sbox_28[41] = 8'd165;
    sbox_28[42] = 8'd229;
    sbox_28[43] = 8'd241;
    sbox_28[44] = 8'd113;
    sbox_28[45] = 8'd216;
    sbox_28[46] = 8'd49;
    sbox_28[47] = 8'd21;
    sbox_28[48] = 8'd4;
    sbox_28[49] = 8'd199;
    sbox_28[50] = 8'd35;
    sbox_28[51] = 8'd195;
    sbox_28[52] = 8'd24;
    sbox_28[53] = 8'd150;
    sbox_28[54] = 8'd5;
    sbox_28[55] = 8'd154;
    sbox_28[56] = 8'd7;
    sbox_28[57] = 8'd18;
    sbox_28[58] = 8'd128;
    sbox_28[59] = 8'd226;
    sbox_28[60] = 8'd235;
    sbox_28[61] = 8'd39;
    sbox_28[62] = 8'd178;
    sbox_28[63] = 8'd117;
    sbox_28[64] = 8'd9;
    sbox_28[65] = 8'd131;
    sbox_28[66] = 8'd44;
    sbox_28[67] = 8'd26;
    sbox_28[68] = 8'd27;
    sbox_28[69] = 8'd110;
    sbox_28[70] = 8'd90;
    sbox_28[71] = 8'd160;
    sbox_28[72] = 8'd82;
    sbox_28[73] = 8'd59;
    sbox_28[74] = 8'd214;
    sbox_28[75] = 8'd179;
    sbox_28[76] = 8'd41;
    sbox_28[77] = 8'd227;
    sbox_28[78] = 8'd47;
    sbox_28[79] = 8'd132;
    sbox_28[80] = 8'd83;
    sbox_28[81] = 8'd209;
    sbox_28[82] = 8'd0;
    sbox_28[83] = 8'd237;
    sbox_28[84] = 8'd32;
    sbox_28[85] = 8'd252;
    sbox_28[86] = 8'd177;
    sbox_28[87] = 8'd91;
    sbox_28[88] = 8'd106;
    sbox_28[89] = 8'd203;
    sbox_28[90] = 8'd190;
    sbox_28[91] = 8'd57;
    sbox_28[92] = 8'd74;
    sbox_28[93] = 8'd76;
    sbox_28[94] = 8'd88;
    sbox_28[95] = 8'd207;
    sbox_28[96] = 8'd208;
    sbox_28[97] = 8'd239;
    sbox_28[98] = 8'd170;
    sbox_28[99] = 8'd251;
    sbox_28[100] = 8'd67;
    sbox_28[101] = 8'd77;
    sbox_28[102] = 8'd51;
    sbox_28[103] = 8'd133;
    sbox_28[104] = 8'd69;
    sbox_28[105] = 8'd249;
    sbox_28[106] = 8'd2;
    sbox_28[107] = 8'd127;
    sbox_28[108] = 8'd80;
    sbox_28[109] = 8'd60;
    sbox_28[110] = 8'd159;
    sbox_28[111] = 8'd168;
    sbox_28[112] = 8'd81;
    sbox_28[113] = 8'd163;
    sbox_28[114] = 8'd64;
    sbox_28[115] = 8'd143;
    sbox_28[116] = 8'd146;
    sbox_28[117] = 8'd157;
    sbox_28[118] = 8'd56;
    sbox_28[119] = 8'd245;
    sbox_28[120] = 8'd188;
    sbox_28[121] = 8'd182;
    sbox_28[122] = 8'd218;
    sbox_28[123] = 8'd33;
    sbox_28[124] = 8'd16;
    sbox_28[125] = 8'd255;
    sbox_28[126] = 8'd243;
    sbox_28[127] = 8'd210;
    sbox_28[128] = 8'd205;
    sbox_28[129] = 8'd12;
    sbox_28[130] = 8'd19;
    sbox_28[131] = 8'd236;
    sbox_28[132] = 8'd95;
    sbox_28[133] = 8'd151;
    sbox_28[134] = 8'd68;
    sbox_28[135] = 8'd23;
    sbox_28[136] = 8'd196;
    sbox_28[137] = 8'd167;
    sbox_28[138] = 8'd126;
    sbox_28[139] = 8'd61;
    sbox_28[140] = 8'd100;
    sbox_28[141] = 8'd93;
    sbox_28[142] = 8'd25;
    sbox_28[143] = 8'd115;
    sbox_28[144] = 8'd96;
    sbox_28[145] = 8'd129;
    sbox_28[146] = 8'd79;
    sbox_28[147] = 8'd220;
    sbox_28[148] = 8'd34;
    sbox_28[149] = 8'd42;
    sbox_28[150] = 8'd144;
    sbox_28[151] = 8'd136;
    sbox_28[152] = 8'd70;
    sbox_28[153] = 8'd238;
    sbox_28[154] = 8'd184;
    sbox_28[155] = 8'd20;
    sbox_28[156] = 8'd222;
    sbox_28[157] = 8'd94;
    sbox_28[158] = 8'd11;
    sbox_28[159] = 8'd219;
    sbox_28[160] = 8'd224;
    sbox_28[161] = 8'd50;
    sbox_28[162] = 8'd58;
    sbox_28[163] = 8'd10;
    sbox_28[164] = 8'd73;
    sbox_28[165] = 8'd6;
    sbox_28[166] = 8'd36;
    sbox_28[167] = 8'd92;
    sbox_28[168] = 8'd194;
    sbox_28[169] = 8'd211;
    sbox_28[170] = 8'd172;
    sbox_28[171] = 8'd98;
    sbox_28[172] = 8'd145;
    sbox_28[173] = 8'd149;
    sbox_28[174] = 8'd228;
    sbox_28[175] = 8'd121;
    sbox_28[176] = 8'd231;
    sbox_28[177] = 8'd200;
    sbox_28[178] = 8'd55;
    sbox_28[179] = 8'd109;
    sbox_28[180] = 8'd141;
    sbox_28[181] = 8'd213;
    sbox_28[182] = 8'd78;
    sbox_28[183] = 8'd169;
    sbox_28[184] = 8'd108;
    sbox_28[185] = 8'd86;
    sbox_28[186] = 8'd244;
    sbox_28[187] = 8'd234;
    sbox_28[188] = 8'd101;
    sbox_28[189] = 8'd122;
    sbox_28[190] = 8'd174;
    sbox_28[191] = 8'd8;
    sbox_28[192] = 8'd186;
    sbox_28[193] = 8'd120;
    sbox_28[194] = 8'd37;
    sbox_28[195] = 8'd46;
    sbox_28[196] = 8'd28;
    sbox_28[197] = 8'd166;
    sbox_28[198] = 8'd180;
    sbox_28[199] = 8'd198;
    sbox_28[200] = 8'd232;
    sbox_28[201] = 8'd221;
    sbox_28[202] = 8'd116;
    sbox_28[203] = 8'd31;
    sbox_28[204] = 8'd75;
    sbox_28[205] = 8'd189;
    sbox_28[206] = 8'd139;
    sbox_28[207] = 8'd138;
    sbox_28[208] = 8'd112;
    sbox_28[209] = 8'd62;
    sbox_28[210] = 8'd181;
    sbox_28[211] = 8'd102;
    sbox_28[212] = 8'd72;
    sbox_28[213] = 8'd3;
    sbox_28[214] = 8'd246;
    sbox_28[215] = 8'd14;
    sbox_28[216] = 8'd97;
    sbox_28[217] = 8'd53;
    sbox_28[218] = 8'd87;
    sbox_28[219] = 8'd185;
    sbox_28[220] = 8'd134;
    sbox_28[221] = 8'd193;
    sbox_28[222] = 8'd29;
    sbox_28[223] = 8'd158;
    sbox_28[224] = 8'd225;
    sbox_28[225] = 8'd248;
    sbox_28[226] = 8'd152;
    sbox_28[227] = 8'd17;
    sbox_28[228] = 8'd105;
    sbox_28[229] = 8'd217;
    sbox_28[230] = 8'd142;
    sbox_28[231] = 8'd148;
    sbox_28[232] = 8'd155;
    sbox_28[233] = 8'd30;
    sbox_28[234] = 8'd135;
    sbox_28[235] = 8'd233;
    sbox_28[236] = 8'd206;
    sbox_28[237] = 8'd85;
    sbox_28[238] = 8'd40;
    sbox_28[239] = 8'd223;
    sbox_28[240] = 8'd140;
    sbox_28[241] = 8'd161;
    sbox_28[242] = 8'd137;
    sbox_28[243] = 8'd13;
    sbox_28[244] = 8'd191;
    sbox_28[245] = 8'd230;
    sbox_28[246] = 8'd66;
    sbox_28[247] = 8'd104;
    sbox_28[248] = 8'd65;
    sbox_28[249] = 8'd153;
    sbox_28[250] = 8'd45;
    sbox_28[251] = 8'd15;
    sbox_28[252] = 8'd176;
    sbox_28[253] = 8'd84;
    sbox_28[254] = 8'd187;
    sbox_28[255] = 8'd22;
    sbox_29[0] = 8'd99;
    sbox_29[1] = 8'd124;
    sbox_29[2] = 8'd119;
    sbox_29[3] = 8'd123;
    sbox_29[4] = 8'd242;
    sbox_29[5] = 8'd107;
    sbox_29[6] = 8'd111;
    sbox_29[7] = 8'd197;
    sbox_29[8] = 8'd48;
    sbox_29[9] = 8'd1;
    sbox_29[10] = 8'd103;
    sbox_29[11] = 8'd43;
    sbox_29[12] = 8'd254;
    sbox_29[13] = 8'd215;
    sbox_29[14] = 8'd171;
    sbox_29[15] = 8'd118;
    sbox_29[16] = 8'd202;
    sbox_29[17] = 8'd130;
    sbox_29[18] = 8'd201;
    sbox_29[19] = 8'd125;
    sbox_29[20] = 8'd250;
    sbox_29[21] = 8'd89;
    sbox_29[22] = 8'd71;
    sbox_29[23] = 8'd240;
    sbox_29[24] = 8'd173;
    sbox_29[25] = 8'd212;
    sbox_29[26] = 8'd162;
    sbox_29[27] = 8'd175;
    sbox_29[28] = 8'd156;
    sbox_29[29] = 8'd164;
    sbox_29[30] = 8'd114;
    sbox_29[31] = 8'd192;
    sbox_29[32] = 8'd183;
    sbox_29[33] = 8'd253;
    sbox_29[34] = 8'd147;
    sbox_29[35] = 8'd38;
    sbox_29[36] = 8'd54;
    sbox_29[37] = 8'd63;
    sbox_29[38] = 8'd247;
    sbox_29[39] = 8'd204;
    sbox_29[40] = 8'd52;
    sbox_29[41] = 8'd165;
    sbox_29[42] = 8'd229;
    sbox_29[43] = 8'd241;
    sbox_29[44] = 8'd113;
    sbox_29[45] = 8'd216;
    sbox_29[46] = 8'd49;
    sbox_29[47] = 8'd21;
    sbox_29[48] = 8'd4;
    sbox_29[49] = 8'd199;
    sbox_29[50] = 8'd35;
    sbox_29[51] = 8'd195;
    sbox_29[52] = 8'd24;
    sbox_29[53] = 8'd150;
    sbox_29[54] = 8'd5;
    sbox_29[55] = 8'd154;
    sbox_29[56] = 8'd7;
    sbox_29[57] = 8'd18;
    sbox_29[58] = 8'd128;
    sbox_29[59] = 8'd226;
    sbox_29[60] = 8'd235;
    sbox_29[61] = 8'd39;
    sbox_29[62] = 8'd178;
    sbox_29[63] = 8'd117;
    sbox_29[64] = 8'd9;
    sbox_29[65] = 8'd131;
    sbox_29[66] = 8'd44;
    sbox_29[67] = 8'd26;
    sbox_29[68] = 8'd27;
    sbox_29[69] = 8'd110;
    sbox_29[70] = 8'd90;
    sbox_29[71] = 8'd160;
    sbox_29[72] = 8'd82;
    sbox_29[73] = 8'd59;
    sbox_29[74] = 8'd214;
    sbox_29[75] = 8'd179;
    sbox_29[76] = 8'd41;
    sbox_29[77] = 8'd227;
    sbox_29[78] = 8'd47;
    sbox_29[79] = 8'd132;
    sbox_29[80] = 8'd83;
    sbox_29[81] = 8'd209;
    sbox_29[82] = 8'd0;
    sbox_29[83] = 8'd237;
    sbox_29[84] = 8'd32;
    sbox_29[85] = 8'd252;
    sbox_29[86] = 8'd177;
    sbox_29[87] = 8'd91;
    sbox_29[88] = 8'd106;
    sbox_29[89] = 8'd203;
    sbox_29[90] = 8'd190;
    sbox_29[91] = 8'd57;
    sbox_29[92] = 8'd74;
    sbox_29[93] = 8'd76;
    sbox_29[94] = 8'd88;
    sbox_29[95] = 8'd207;
    sbox_29[96] = 8'd208;
    sbox_29[97] = 8'd239;
    sbox_29[98] = 8'd170;
    sbox_29[99] = 8'd251;
    sbox_29[100] = 8'd67;
    sbox_29[101] = 8'd77;
    sbox_29[102] = 8'd51;
    sbox_29[103] = 8'd133;
    sbox_29[104] = 8'd69;
    sbox_29[105] = 8'd249;
    sbox_29[106] = 8'd2;
    sbox_29[107] = 8'd127;
    sbox_29[108] = 8'd80;
    sbox_29[109] = 8'd60;
    sbox_29[110] = 8'd159;
    sbox_29[111] = 8'd168;
    sbox_29[112] = 8'd81;
    sbox_29[113] = 8'd163;
    sbox_29[114] = 8'd64;
    sbox_29[115] = 8'd143;
    sbox_29[116] = 8'd146;
    sbox_29[117] = 8'd157;
    sbox_29[118] = 8'd56;
    sbox_29[119] = 8'd245;
    sbox_29[120] = 8'd188;
    sbox_29[121] = 8'd182;
    sbox_29[122] = 8'd218;
    sbox_29[123] = 8'd33;
    sbox_29[124] = 8'd16;
    sbox_29[125] = 8'd255;
    sbox_29[126] = 8'd243;
    sbox_29[127] = 8'd210;
    sbox_29[128] = 8'd205;
    sbox_29[129] = 8'd12;
    sbox_29[130] = 8'd19;
    sbox_29[131] = 8'd236;
    sbox_29[132] = 8'd95;
    sbox_29[133] = 8'd151;
    sbox_29[134] = 8'd68;
    sbox_29[135] = 8'd23;
    sbox_29[136] = 8'd196;
    sbox_29[137] = 8'd167;
    sbox_29[138] = 8'd126;
    sbox_29[139] = 8'd61;
    sbox_29[140] = 8'd100;
    sbox_29[141] = 8'd93;
    sbox_29[142] = 8'd25;
    sbox_29[143] = 8'd115;
    sbox_29[144] = 8'd96;
    sbox_29[145] = 8'd129;
    sbox_29[146] = 8'd79;
    sbox_29[147] = 8'd220;
    sbox_29[148] = 8'd34;
    sbox_29[149] = 8'd42;
    sbox_29[150] = 8'd144;
    sbox_29[151] = 8'd136;
    sbox_29[152] = 8'd70;
    sbox_29[153] = 8'd238;
    sbox_29[154] = 8'd184;
    sbox_29[155] = 8'd20;
    sbox_29[156] = 8'd222;
    sbox_29[157] = 8'd94;
    sbox_29[158] = 8'd11;
    sbox_29[159] = 8'd219;
    sbox_29[160] = 8'd224;
    sbox_29[161] = 8'd50;
    sbox_29[162] = 8'd58;
    sbox_29[163] = 8'd10;
    sbox_29[164] = 8'd73;
    sbox_29[165] = 8'd6;
    sbox_29[166] = 8'd36;
    sbox_29[167] = 8'd92;
    sbox_29[168] = 8'd194;
    sbox_29[169] = 8'd211;
    sbox_29[170] = 8'd172;
    sbox_29[171] = 8'd98;
    sbox_29[172] = 8'd145;
    sbox_29[173] = 8'd149;
    sbox_29[174] = 8'd228;
    sbox_29[175] = 8'd121;
    sbox_29[176] = 8'd231;
    sbox_29[177] = 8'd200;
    sbox_29[178] = 8'd55;
    sbox_29[179] = 8'd109;
    sbox_29[180] = 8'd141;
    sbox_29[181] = 8'd213;
    sbox_29[182] = 8'd78;
    sbox_29[183] = 8'd169;
    sbox_29[184] = 8'd108;
    sbox_29[185] = 8'd86;
    sbox_29[186] = 8'd244;
    sbox_29[187] = 8'd234;
    sbox_29[188] = 8'd101;
    sbox_29[189] = 8'd122;
    sbox_29[190] = 8'd174;
    sbox_29[191] = 8'd8;
    sbox_29[192] = 8'd186;
    sbox_29[193] = 8'd120;
    sbox_29[194] = 8'd37;
    sbox_29[195] = 8'd46;
    sbox_29[196] = 8'd28;
    sbox_29[197] = 8'd166;
    sbox_29[198] = 8'd180;
    sbox_29[199] = 8'd198;
    sbox_29[200] = 8'd232;
    sbox_29[201] = 8'd221;
    sbox_29[202] = 8'd116;
    sbox_29[203] = 8'd31;
    sbox_29[204] = 8'd75;
    sbox_29[205] = 8'd189;
    sbox_29[206] = 8'd139;
    sbox_29[207] = 8'd138;
    sbox_29[208] = 8'd112;
    sbox_29[209] = 8'd62;
    sbox_29[210] = 8'd181;
    sbox_29[211] = 8'd102;
    sbox_29[212] = 8'd72;
    sbox_29[213] = 8'd3;
    sbox_29[214] = 8'd246;
    sbox_29[215] = 8'd14;
    sbox_29[216] = 8'd97;
    sbox_29[217] = 8'd53;
    sbox_29[218] = 8'd87;
    sbox_29[219] = 8'd185;
    sbox_29[220] = 8'd134;
    sbox_29[221] = 8'd193;
    sbox_29[222] = 8'd29;
    sbox_29[223] = 8'd158;
    sbox_29[224] = 8'd225;
    sbox_29[225] = 8'd248;
    sbox_29[226] = 8'd152;
    sbox_29[227] = 8'd17;
    sbox_29[228] = 8'd105;
    sbox_29[229] = 8'd217;
    sbox_29[230] = 8'd142;
    sbox_29[231] = 8'd148;
    sbox_29[232] = 8'd155;
    sbox_29[233] = 8'd30;
    sbox_29[234] = 8'd135;
    sbox_29[235] = 8'd233;
    sbox_29[236] = 8'd206;
    sbox_29[237] = 8'd85;
    sbox_29[238] = 8'd40;
    sbox_29[239] = 8'd223;
    sbox_29[240] = 8'd140;
    sbox_29[241] = 8'd161;
    sbox_29[242] = 8'd137;
    sbox_29[243] = 8'd13;
    sbox_29[244] = 8'd191;
    sbox_29[245] = 8'd230;
    sbox_29[246] = 8'd66;
    sbox_29[247] = 8'd104;
    sbox_29[248] = 8'd65;
    sbox_29[249] = 8'd153;
    sbox_29[250] = 8'd45;
    sbox_29[251] = 8'd15;
    sbox_29[252] = 8'd176;
    sbox_29[253] = 8'd84;
    sbox_29[254] = 8'd187;
    sbox_29[255] = 8'd22;
    sbox_30[0] = 8'd99;
    sbox_30[1] = 8'd124;
    sbox_30[2] = 8'd119;
    sbox_30[3] = 8'd123;
    sbox_30[4] = 8'd242;
    sbox_30[5] = 8'd107;
    sbox_30[6] = 8'd111;
    sbox_30[7] = 8'd197;
    sbox_30[8] = 8'd48;
    sbox_30[9] = 8'd1;
    sbox_30[10] = 8'd103;
    sbox_30[11] = 8'd43;
    sbox_30[12] = 8'd254;
    sbox_30[13] = 8'd215;
    sbox_30[14] = 8'd171;
    sbox_30[15] = 8'd118;
    sbox_30[16] = 8'd202;
    sbox_30[17] = 8'd130;
    sbox_30[18] = 8'd201;
    sbox_30[19] = 8'd125;
    sbox_30[20] = 8'd250;
    sbox_30[21] = 8'd89;
    sbox_30[22] = 8'd71;
    sbox_30[23] = 8'd240;
    sbox_30[24] = 8'd173;
    sbox_30[25] = 8'd212;
    sbox_30[26] = 8'd162;
    sbox_30[27] = 8'd175;
    sbox_30[28] = 8'd156;
    sbox_30[29] = 8'd164;
    sbox_30[30] = 8'd114;
    sbox_30[31] = 8'd192;
    sbox_30[32] = 8'd183;
    sbox_30[33] = 8'd253;
    sbox_30[34] = 8'd147;
    sbox_30[35] = 8'd38;
    sbox_30[36] = 8'd54;
    sbox_30[37] = 8'd63;
    sbox_30[38] = 8'd247;
    sbox_30[39] = 8'd204;
    sbox_30[40] = 8'd52;
    sbox_30[41] = 8'd165;
    sbox_30[42] = 8'd229;
    sbox_30[43] = 8'd241;
    sbox_30[44] = 8'd113;
    sbox_30[45] = 8'd216;
    sbox_30[46] = 8'd49;
    sbox_30[47] = 8'd21;
    sbox_30[48] = 8'd4;
    sbox_30[49] = 8'd199;
    sbox_30[50] = 8'd35;
    sbox_30[51] = 8'd195;
    sbox_30[52] = 8'd24;
    sbox_30[53] = 8'd150;
    sbox_30[54] = 8'd5;
    sbox_30[55] = 8'd154;
    sbox_30[56] = 8'd7;
    sbox_30[57] = 8'd18;
    sbox_30[58] = 8'd128;
    sbox_30[59] = 8'd226;
    sbox_30[60] = 8'd235;
    sbox_30[61] = 8'd39;
    sbox_30[62] = 8'd178;
    sbox_30[63] = 8'd117;
    sbox_30[64] = 8'd9;
    sbox_30[65] = 8'd131;
    sbox_30[66] = 8'd44;
    sbox_30[67] = 8'd26;
    sbox_30[68] = 8'd27;
    sbox_30[69] = 8'd110;
    sbox_30[70] = 8'd90;
    sbox_30[71] = 8'd160;
    sbox_30[72] = 8'd82;
    sbox_30[73] = 8'd59;
    sbox_30[74] = 8'd214;
    sbox_30[75] = 8'd179;
    sbox_30[76] = 8'd41;
    sbox_30[77] = 8'd227;
    sbox_30[78] = 8'd47;
    sbox_30[79] = 8'd132;
    sbox_30[80] = 8'd83;
    sbox_30[81] = 8'd209;
    sbox_30[82] = 8'd0;
    sbox_30[83] = 8'd237;
    sbox_30[84] = 8'd32;
    sbox_30[85] = 8'd252;
    sbox_30[86] = 8'd177;
    sbox_30[87] = 8'd91;
    sbox_30[88] = 8'd106;
    sbox_30[89] = 8'd203;
    sbox_30[90] = 8'd190;
    sbox_30[91] = 8'd57;
    sbox_30[92] = 8'd74;
    sbox_30[93] = 8'd76;
    sbox_30[94] = 8'd88;
    sbox_30[95] = 8'd207;
    sbox_30[96] = 8'd208;
    sbox_30[97] = 8'd239;
    sbox_30[98] = 8'd170;
    sbox_30[99] = 8'd251;
    sbox_30[100] = 8'd67;
    sbox_30[101] = 8'd77;
    sbox_30[102] = 8'd51;
    sbox_30[103] = 8'd133;
    sbox_30[104] = 8'd69;
    sbox_30[105] = 8'd249;
    sbox_30[106] = 8'd2;
    sbox_30[107] = 8'd127;
    sbox_30[108] = 8'd80;
    sbox_30[109] = 8'd60;
    sbox_30[110] = 8'd159;
    sbox_30[111] = 8'd168;
    sbox_30[112] = 8'd81;
    sbox_30[113] = 8'd163;
    sbox_30[114] = 8'd64;
    sbox_30[115] = 8'd143;
    sbox_30[116] = 8'd146;
    sbox_30[117] = 8'd157;
    sbox_30[118] = 8'd56;
    sbox_30[119] = 8'd245;
    sbox_30[120] = 8'd188;
    sbox_30[121] = 8'd182;
    sbox_30[122] = 8'd218;
    sbox_30[123] = 8'd33;
    sbox_30[124] = 8'd16;
    sbox_30[125] = 8'd255;
    sbox_30[126] = 8'd243;
    sbox_30[127] = 8'd210;
    sbox_30[128] = 8'd205;
    sbox_30[129] = 8'd12;
    sbox_30[130] = 8'd19;
    sbox_30[131] = 8'd236;
    sbox_30[132] = 8'd95;
    sbox_30[133] = 8'd151;
    sbox_30[134] = 8'd68;
    sbox_30[135] = 8'd23;
    sbox_30[136] = 8'd196;
    sbox_30[137] = 8'd167;
    sbox_30[138] = 8'd126;
    sbox_30[139] = 8'd61;
    sbox_30[140] = 8'd100;
    sbox_30[141] = 8'd93;
    sbox_30[142] = 8'd25;
    sbox_30[143] = 8'd115;
    sbox_30[144] = 8'd96;
    sbox_30[145] = 8'd129;
    sbox_30[146] = 8'd79;
    sbox_30[147] = 8'd220;
    sbox_30[148] = 8'd34;
    sbox_30[149] = 8'd42;
    sbox_30[150] = 8'd144;
    sbox_30[151] = 8'd136;
    sbox_30[152] = 8'd70;
    sbox_30[153] = 8'd238;
    sbox_30[154] = 8'd184;
    sbox_30[155] = 8'd20;
    sbox_30[156] = 8'd222;
    sbox_30[157] = 8'd94;
    sbox_30[158] = 8'd11;
    sbox_30[159] = 8'd219;
    sbox_30[160] = 8'd224;
    sbox_30[161] = 8'd50;
    sbox_30[162] = 8'd58;
    sbox_30[163] = 8'd10;
    sbox_30[164] = 8'd73;
    sbox_30[165] = 8'd6;
    sbox_30[166] = 8'd36;
    sbox_30[167] = 8'd92;
    sbox_30[168] = 8'd194;
    sbox_30[169] = 8'd211;
    sbox_30[170] = 8'd172;
    sbox_30[171] = 8'd98;
    sbox_30[172] = 8'd145;
    sbox_30[173] = 8'd149;
    sbox_30[174] = 8'd228;
    sbox_30[175] = 8'd121;
    sbox_30[176] = 8'd231;
    sbox_30[177] = 8'd200;
    sbox_30[178] = 8'd55;
    sbox_30[179] = 8'd109;
    sbox_30[180] = 8'd141;
    sbox_30[181] = 8'd213;
    sbox_30[182] = 8'd78;
    sbox_30[183] = 8'd169;
    sbox_30[184] = 8'd108;
    sbox_30[185] = 8'd86;
    sbox_30[186] = 8'd244;
    sbox_30[187] = 8'd234;
    sbox_30[188] = 8'd101;
    sbox_30[189] = 8'd122;
    sbox_30[190] = 8'd174;
    sbox_30[191] = 8'd8;
    sbox_30[192] = 8'd186;
    sbox_30[193] = 8'd120;
    sbox_30[194] = 8'd37;
    sbox_30[195] = 8'd46;
    sbox_30[196] = 8'd28;
    sbox_30[197] = 8'd166;
    sbox_30[198] = 8'd180;
    sbox_30[199] = 8'd198;
    sbox_30[200] = 8'd232;
    sbox_30[201] = 8'd221;
    sbox_30[202] = 8'd116;
    sbox_30[203] = 8'd31;
    sbox_30[204] = 8'd75;
    sbox_30[205] = 8'd189;
    sbox_30[206] = 8'd139;
    sbox_30[207] = 8'd138;
    sbox_30[208] = 8'd112;
    sbox_30[209] = 8'd62;
    sbox_30[210] = 8'd181;
    sbox_30[211] = 8'd102;
    sbox_30[212] = 8'd72;
    sbox_30[213] = 8'd3;
    sbox_30[214] = 8'd246;
    sbox_30[215] = 8'd14;
    sbox_30[216] = 8'd97;
    sbox_30[217] = 8'd53;
    sbox_30[218] = 8'd87;
    sbox_30[219] = 8'd185;
    sbox_30[220] = 8'd134;
    sbox_30[221] = 8'd193;
    sbox_30[222] = 8'd29;
    sbox_30[223] = 8'd158;
    sbox_30[224] = 8'd225;
    sbox_30[225] = 8'd248;
    sbox_30[226] = 8'd152;
    sbox_30[227] = 8'd17;
    sbox_30[228] = 8'd105;
    sbox_30[229] = 8'd217;
    sbox_30[230] = 8'd142;
    sbox_30[231] = 8'd148;
    sbox_30[232] = 8'd155;
    sbox_30[233] = 8'd30;
    sbox_30[234] = 8'd135;
    sbox_30[235] = 8'd233;
    sbox_30[236] = 8'd206;
    sbox_30[237] = 8'd85;
    sbox_30[238] = 8'd40;
    sbox_30[239] = 8'd223;
    sbox_30[240] = 8'd140;
    sbox_30[241] = 8'd161;
    sbox_30[242] = 8'd137;
    sbox_30[243] = 8'd13;
    sbox_30[244] = 8'd191;
    sbox_30[245] = 8'd230;
    sbox_30[246] = 8'd66;
    sbox_30[247] = 8'd104;
    sbox_30[248] = 8'd65;
    sbox_30[249] = 8'd153;
    sbox_30[250] = 8'd45;
    sbox_30[251] = 8'd15;
    sbox_30[252] = 8'd176;
    sbox_30[253] = 8'd84;
    sbox_30[254] = 8'd187;
    sbox_30[255] = 8'd22;
    sbox_31[0] = 8'd99;
    sbox_31[1] = 8'd124;
    sbox_31[2] = 8'd119;
    sbox_31[3] = 8'd123;
    sbox_31[4] = 8'd242;
    sbox_31[5] = 8'd107;
    sbox_31[6] = 8'd111;
    sbox_31[7] = 8'd197;
    sbox_31[8] = 8'd48;
    sbox_31[9] = 8'd1;
    sbox_31[10] = 8'd103;
    sbox_31[11] = 8'd43;
    sbox_31[12] = 8'd254;
    sbox_31[13] = 8'd215;
    sbox_31[14] = 8'd171;
    sbox_31[15] = 8'd118;
    sbox_31[16] = 8'd202;
    sbox_31[17] = 8'd130;
    sbox_31[18] = 8'd201;
    sbox_31[19] = 8'd125;
    sbox_31[20] = 8'd250;
    sbox_31[21] = 8'd89;
    sbox_31[22] = 8'd71;
    sbox_31[23] = 8'd240;
    sbox_31[24] = 8'd173;
    sbox_31[25] = 8'd212;
    sbox_31[26] = 8'd162;
    sbox_31[27] = 8'd175;
    sbox_31[28] = 8'd156;
    sbox_31[29] = 8'd164;
    sbox_31[30] = 8'd114;
    sbox_31[31] = 8'd192;
    sbox_31[32] = 8'd183;
    sbox_31[33] = 8'd253;
    sbox_31[34] = 8'd147;
    sbox_31[35] = 8'd38;
    sbox_31[36] = 8'd54;
    sbox_31[37] = 8'd63;
    sbox_31[38] = 8'd247;
    sbox_31[39] = 8'd204;
    sbox_31[40] = 8'd52;
    sbox_31[41] = 8'd165;
    sbox_31[42] = 8'd229;
    sbox_31[43] = 8'd241;
    sbox_31[44] = 8'd113;
    sbox_31[45] = 8'd216;
    sbox_31[46] = 8'd49;
    sbox_31[47] = 8'd21;
    sbox_31[48] = 8'd4;
    sbox_31[49] = 8'd199;
    sbox_31[50] = 8'd35;
    sbox_31[51] = 8'd195;
    sbox_31[52] = 8'd24;
    sbox_31[53] = 8'd150;
    sbox_31[54] = 8'd5;
    sbox_31[55] = 8'd154;
    sbox_31[56] = 8'd7;
    sbox_31[57] = 8'd18;
    sbox_31[58] = 8'd128;
    sbox_31[59] = 8'd226;
    sbox_31[60] = 8'd235;
    sbox_31[61] = 8'd39;
    sbox_31[62] = 8'd178;
    sbox_31[63] = 8'd117;
    sbox_31[64] = 8'd9;
    sbox_31[65] = 8'd131;
    sbox_31[66] = 8'd44;
    sbox_31[67] = 8'd26;
    sbox_31[68] = 8'd27;
    sbox_31[69] = 8'd110;
    sbox_31[70] = 8'd90;
    sbox_31[71] = 8'd160;
    sbox_31[72] = 8'd82;
    sbox_31[73] = 8'd59;
    sbox_31[74] = 8'd214;
    sbox_31[75] = 8'd179;
    sbox_31[76] = 8'd41;
    sbox_31[77] = 8'd227;
    sbox_31[78] = 8'd47;
    sbox_31[79] = 8'd132;
    sbox_31[80] = 8'd83;
    sbox_31[81] = 8'd209;
    sbox_31[82] = 8'd0;
    sbox_31[83] = 8'd237;
    sbox_31[84] = 8'd32;
    sbox_31[85] = 8'd252;
    sbox_31[86] = 8'd177;
    sbox_31[87] = 8'd91;
    sbox_31[88] = 8'd106;
    sbox_31[89] = 8'd203;
    sbox_31[90] = 8'd190;
    sbox_31[91] = 8'd57;
    sbox_31[92] = 8'd74;
    sbox_31[93] = 8'd76;
    sbox_31[94] = 8'd88;
    sbox_31[95] = 8'd207;
    sbox_31[96] = 8'd208;
    sbox_31[97] = 8'd239;
    sbox_31[98] = 8'd170;
    sbox_31[99] = 8'd251;
    sbox_31[100] = 8'd67;
    sbox_31[101] = 8'd77;
    sbox_31[102] = 8'd51;
    sbox_31[103] = 8'd133;
    sbox_31[104] = 8'd69;
    sbox_31[105] = 8'd249;
    sbox_31[106] = 8'd2;
    sbox_31[107] = 8'd127;
    sbox_31[108] = 8'd80;
    sbox_31[109] = 8'd60;
    sbox_31[110] = 8'd159;
    sbox_31[111] = 8'd168;
    sbox_31[112] = 8'd81;
    sbox_31[113] = 8'd163;
    sbox_31[114] = 8'd64;
    sbox_31[115] = 8'd143;
    sbox_31[116] = 8'd146;
    sbox_31[117] = 8'd157;
    sbox_31[118] = 8'd56;
    sbox_31[119] = 8'd245;
    sbox_31[120] = 8'd188;
    sbox_31[121] = 8'd182;
    sbox_31[122] = 8'd218;
    sbox_31[123] = 8'd33;
    sbox_31[124] = 8'd16;
    sbox_31[125] = 8'd255;
    sbox_31[126] = 8'd243;
    sbox_31[127] = 8'd210;
    sbox_31[128] = 8'd205;
    sbox_31[129] = 8'd12;
    sbox_31[130] = 8'd19;
    sbox_31[131] = 8'd236;
    sbox_31[132] = 8'd95;
    sbox_31[133] = 8'd151;
    sbox_31[134] = 8'd68;
    sbox_31[135] = 8'd23;
    sbox_31[136] = 8'd196;
    sbox_31[137] = 8'd167;
    sbox_31[138] = 8'd126;
    sbox_31[139] = 8'd61;
    sbox_31[140] = 8'd100;
    sbox_31[141] = 8'd93;
    sbox_31[142] = 8'd25;
    sbox_31[143] = 8'd115;
    sbox_31[144] = 8'd96;
    sbox_31[145] = 8'd129;
    sbox_31[146] = 8'd79;
    sbox_31[147] = 8'd220;
    sbox_31[148] = 8'd34;
    sbox_31[149] = 8'd42;
    sbox_31[150] = 8'd144;
    sbox_31[151] = 8'd136;
    sbox_31[152] = 8'd70;
    sbox_31[153] = 8'd238;
    sbox_31[154] = 8'd184;
    sbox_31[155] = 8'd20;
    sbox_31[156] = 8'd222;
    sbox_31[157] = 8'd94;
    sbox_31[158] = 8'd11;
    sbox_31[159] = 8'd219;
    sbox_31[160] = 8'd224;
    sbox_31[161] = 8'd50;
    sbox_31[162] = 8'd58;
    sbox_31[163] = 8'd10;
    sbox_31[164] = 8'd73;
    sbox_31[165] = 8'd6;
    sbox_31[166] = 8'd36;
    sbox_31[167] = 8'd92;
    sbox_31[168] = 8'd194;
    sbox_31[169] = 8'd211;
    sbox_31[170] = 8'd172;
    sbox_31[171] = 8'd98;
    sbox_31[172] = 8'd145;
    sbox_31[173] = 8'd149;
    sbox_31[174] = 8'd228;
    sbox_31[175] = 8'd121;
    sbox_31[176] = 8'd231;
    sbox_31[177] = 8'd200;
    sbox_31[178] = 8'd55;
    sbox_31[179] = 8'd109;
    sbox_31[180] = 8'd141;
    sbox_31[181] = 8'd213;
    sbox_31[182] = 8'd78;
    sbox_31[183] = 8'd169;
    sbox_31[184] = 8'd108;
    sbox_31[185] = 8'd86;
    sbox_31[186] = 8'd244;
    sbox_31[187] = 8'd234;
    sbox_31[188] = 8'd101;
    sbox_31[189] = 8'd122;
    sbox_31[190] = 8'd174;
    sbox_31[191] = 8'd8;
    sbox_31[192] = 8'd186;
    sbox_31[193] = 8'd120;
    sbox_31[194] = 8'd37;
    sbox_31[195] = 8'd46;
    sbox_31[196] = 8'd28;
    sbox_31[197] = 8'd166;
    sbox_31[198] = 8'd180;
    sbox_31[199] = 8'd198;
    sbox_31[200] = 8'd232;
    sbox_31[201] = 8'd221;
    sbox_31[202] = 8'd116;
    sbox_31[203] = 8'd31;
    sbox_31[204] = 8'd75;
    sbox_31[205] = 8'd189;
    sbox_31[206] = 8'd139;
    sbox_31[207] = 8'd138;
    sbox_31[208] = 8'd112;
    sbox_31[209] = 8'd62;
    sbox_31[210] = 8'd181;
    sbox_31[211] = 8'd102;
    sbox_31[212] = 8'd72;
    sbox_31[213] = 8'd3;
    sbox_31[214] = 8'd246;
    sbox_31[215] = 8'd14;
    sbox_31[216] = 8'd97;
    sbox_31[217] = 8'd53;
    sbox_31[218] = 8'd87;
    sbox_31[219] = 8'd185;
    sbox_31[220] = 8'd134;
    sbox_31[221] = 8'd193;
    sbox_31[222] = 8'd29;
    sbox_31[223] = 8'd158;
    sbox_31[224] = 8'd225;
    sbox_31[225] = 8'd248;
    sbox_31[226] = 8'd152;
    sbox_31[227] = 8'd17;
    sbox_31[228] = 8'd105;
    sbox_31[229] = 8'd217;
    sbox_31[230] = 8'd142;
    sbox_31[231] = 8'd148;
    sbox_31[232] = 8'd155;
    sbox_31[233] = 8'd30;
    sbox_31[234] = 8'd135;
    sbox_31[235] = 8'd233;
    sbox_31[236] = 8'd206;
    sbox_31[237] = 8'd85;
    sbox_31[238] = 8'd40;
    sbox_31[239] = 8'd223;
    sbox_31[240] = 8'd140;
    sbox_31[241] = 8'd161;
    sbox_31[242] = 8'd137;
    sbox_31[243] = 8'd13;
    sbox_31[244] = 8'd191;
    sbox_31[245] = 8'd230;
    sbox_31[246] = 8'd66;
    sbox_31[247] = 8'd104;
    sbox_31[248] = 8'd65;
    sbox_31[249] = 8'd153;
    sbox_31[250] = 8'd45;
    sbox_31[251] = 8'd15;
    sbox_31[252] = 8'd176;
    sbox_31[253] = 8'd84;
    sbox_31[254] = 8'd187;
    sbox_31[255] = 8'd22;
end
    assign lookup_sbox_0_enable = (1'd0);
    assign lookup_sbox_0_0 = (1'd0);
    assign lookup_sbox_1_enable = (1'd0);
    assign lookup_sbox_1_0 = (1'd0);
    assign lookup_sbox_2_enable = (1'd0);
    assign lookup_sbox_2_0 = (1'd0);
    assign lookup_sbox_3_enable = (1'd0);
    assign lookup_sbox_3_0 = (1'd0);
    assign lookup_sbox_4_enable = (1'd0);
    assign lookup_sbox_4_0 = (1'd0);
    assign lookup_sbox_5_enable = (1'd0);
    assign lookup_sbox_5_0 = (1'd0);
    assign lookup_sbox_6_enable = (1'd0);
    assign lookup_sbox_6_0 = (1'd0);
    assign lookup_sbox_7_enable = (1'd0);
    assign lookup_sbox_7_0 = (1'd0);
    assign lookup_sbox_8_enable = (1'd0);
    assign lookup_sbox_8_0 = (1'd0);
    assign lookup_sbox_9_enable = (1'd0);
    assign lookup_sbox_9_0 = (1'd0);
    assign lookup_sbox_10_enable = (1'd0);
    assign lookup_sbox_10_0 = (1'd0);
    assign lookup_sbox_11_enable = (1'd0);
    assign lookup_sbox_11_0 = (1'd0);
    assign lookup_sbox_12_enable = (1'd0);
    assign lookup_sbox_12_0 = (1'd0);
    assign lookup_sbox_13_enable = ((control_194_37)||(1'd0));
    assign lookup_sbox_13_0 = ((control_194_37)?({(operation_194_3046[7:0])}):(1'd0));
    assign lookup_sbox_14_enable = ((control_194_10)||((control_194_37)||(1'd0)));
    assign lookup_sbox_14_0 = ((control_194_10)?({(operation_194_1759[7:0])}):((control_194_37)?({(operation_194_3044[7:0])}):(1'd0)));
    assign lookup_sbox_15_enable = ((control_194_10)||((control_194_37)||(1'd0)));
    assign lookup_sbox_15_0 = ((control_194_10)?({(operation_194_1757[7:0])}):((control_194_37)?({(operation_194_3042[7:0])}):(1'd0)));
    assign lookup_sbox_16_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_16_0 = ((control_194_1)?({(operation_194_127[7:0])}):((control_194_10)?({(operation_194_1755[7:0])}):((control_194_19)?({(operation_194_2188[7:0])}):((control_194_28)?({(operation_194_2617[7:0])}):((control_194_37)?({(operation_194_3040[7:0])}):((control_194_46)?({(operation_194_3475[7:0])}):((control_194_55)?({(operation_194_3904[7:0])}):((control_194_64)?({(operation_194_4333[7:0])}):((control_194_73)?({(operation_194_4762[7:0])}):((control_194_82)?({(operation_194_5191[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_17_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_17_0 = ((control_194_1)?({(operation_194_111[7:0])}):((control_194_10)?({(operation_194_1753[7:0])}):((control_194_19)?({(operation_194_2186[7:0])}):((control_194_28)?({(operation_194_2615[7:0])}):((control_194_37)?({(operation_194_3038[7:0])}):((control_194_46)?({(operation_194_3473[7:0])}):((control_194_55)?({(operation_194_3902[7:0])}):((control_194_64)?({(operation_194_4331[7:0])}):((control_194_73)?({(operation_194_4760[7:0])}):((control_194_82)?({(operation_194_5189[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_18_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_18_0 = ((control_194_1)?({(operation_194_95[7:0])}):((control_194_10)?({(operation_194_1751[7:0])}):((control_194_19)?({(operation_194_2184[7:0])}):((control_194_28)?({(operation_194_2613[7:0])}):((control_194_37)?({(operation_194_3036[7:0])}):((control_194_46)?({(operation_194_3471[7:0])}):((control_194_55)?({(operation_194_3900[7:0])}):((control_194_64)?({(operation_194_4329[7:0])}):((control_194_73)?({(operation_194_4758[7:0])}):((control_194_82)?({(operation_194_5187[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_19_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_19_0 = ((control_194_1)?({(operation_194_79[7:0])}):((control_194_10)?({(operation_194_1749[7:0])}):((control_194_19)?({(operation_194_2182[7:0])}):((control_194_28)?({(operation_194_2611[7:0])}):((control_194_37)?({(operation_194_3034[7:0])}):((control_194_46)?({(operation_194_3469[7:0])}):((control_194_55)?({(operation_194_3898[7:0])}):((control_194_64)?({(operation_194_4327[7:0])}):((control_194_73)?({(operation_194_4756[7:0])}):((control_194_82)?({(operation_194_5185[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_20_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_20_0 = ((control_194_1)?({(operation_194_63[7:0])}):((control_194_10)?({(operation_194_1747[7:0])}):((control_194_19)?({(operation_194_2180[7:0])}):((control_194_28)?({(operation_194_2609[7:0])}):((control_194_37)?({(operation_194_3032[7:0])}):((control_194_46)?({(operation_194_3467[7:0])}):((control_194_55)?({(operation_194_3896[7:0])}):((control_194_64)?({(operation_194_4325[7:0])}):((control_194_73)?({(operation_194_4754[7:0])}):((control_194_82)?({(operation_194_5183[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_21_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_21_0 = ((control_194_1)?({(operation_194_47[7:0])}):((control_194_10)?({(operation_194_1745[7:0])}):((control_194_19)?({(operation_194_2178[7:0])}):((control_194_28)?({(operation_194_2607[7:0])}):((control_194_37)?({(operation_194_2992[7:0])}):((control_194_46)?({(operation_194_3465[7:0])}):((control_194_55)?({(operation_194_3894[7:0])}):((control_194_64)?({(operation_194_4323[7:0])}):((control_194_73)?({(operation_194_4752[7:0])}):((control_194_82)?({(operation_194_5181[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_22_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_22_0 = ((control_194_1)?({(operation_194_31[7:0])}):((control_194_10)?({(operation_194_1705[7:0])}):((control_194_19)?({(operation_194_2176[7:0])}):((control_194_28)?({(operation_194_2605[7:0])}):((control_194_37)?({(operation_194_2994[7:0])}):((control_194_46)?({(operation_194_3463[7:0])}):((control_194_55)?({(operation_194_3892[7:0])}):((control_194_64)?({(operation_194_4321[7:0])}):((control_194_73)?({(operation_194_4750[7:0])}):((control_194_82)?({(operation_194_5179[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_23_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_23_0 = ((control_194_1)?({(operation_194_15[7:0])}):((control_194_10)?({(operation_194_1707[7:0])}):((control_194_19)?({(operation_194_2174[7:0])}):((control_194_28)?({(operation_194_2603[7:0])}):((control_194_37)?({(operation_194_2996[7:0])}):((control_194_46)?({(operation_194_3461[7:0])}):((control_194_55)?({(operation_194_3890[7:0])}):((control_194_64)?({(operation_194_4319[7:0])}):((control_194_73)?({(operation_194_4748[7:0])}):((control_194_82)?({(operation_194_5177[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_24_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_24_0 = ((control_194_1)?({(operation_194_7[7:0])}):((control_194_10)?({(operation_194_1709[7:0])}):((control_194_19)?({(operation_194_2134[7:0])}):((control_194_28)?({(operation_194_2563[7:0])}):((control_194_37)?({(operation_194_2998[7:0])}):((control_194_46)?({(operation_194_3421[7:0])}):((control_194_55)?({(operation_194_3850[7:0])}):((control_194_64)?({(operation_194_4279[7:0])}):((control_194_73)?({(operation_194_4708[7:0])}):((control_194_82)?({(operation_194_5137[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_25_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_25_0 = ((control_194_1)?({(operation_194_23[7:0])}):((control_194_10)?({(operation_194_1711[7:0])}):((control_194_19)?({(operation_194_2136[7:0])}):((control_194_28)?({(operation_194_2565[7:0])}):((control_194_37)?({(operation_194_3000[7:0])}):((control_194_46)?({(operation_194_3423[7:0])}):((control_194_55)?({(operation_194_3852[7:0])}):((control_194_64)?({(operation_194_4281[7:0])}):((control_194_73)?({(operation_194_4710[7:0])}):((control_194_82)?({(operation_194_5139[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_26_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_26_0 = ((control_194_1)?({(operation_194_39[7:0])}):((control_194_10)?({(operation_194_1713[7:0])}):((control_194_19)?({(operation_194_2138[7:0])}):((control_194_28)?({(operation_194_2567[7:0])}):((control_194_37)?({(operation_194_3002[7:0])}):((control_194_46)?({(operation_194_3425[7:0])}):((control_194_55)?({(operation_194_3854[7:0])}):((control_194_64)?({(operation_194_4283[7:0])}):((control_194_73)?({(operation_194_4712[7:0])}):((control_194_82)?({(operation_194_5141[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_27_enable = ((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_73)||((control_194_82)||(1'd0)))))))))));
    assign lookup_sbox_27_0 = ((control_194_1)?({(operation_194_55[7:0])}):((control_194_10)?({(operation_194_1715[7:0])}):((control_194_19)?({(operation_194_2140[7:0])}):((control_194_28)?({(operation_194_2569[7:0])}):((control_194_37)?({(operation_194_2986[7:0])}):((control_194_46)?({(operation_194_3427[7:0])}):((control_194_55)?({(operation_194_3856[7:0])}):((control_194_64)?({(operation_194_4285[7:0])}):((control_194_73)?({(operation_194_4714[7:0])}):((control_194_82)?({(operation_194_5143[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_28_enable = ((control_194_0)||((control_194_1)||((control_194_10)||((control_194_19)||((control_194_28)||((control_194_21)||((control_194_37)||((control_194_46)||((control_194_55)||((control_194_64)||((control_194_42)||((control_194_73)||((control_194_82)||(1'd0))))))))))))));
    assign lookup_sbox_28_0 = ((control_194_0)?({(operation_194_124[103:96])}):((control_194_1)?({(operation_194_71[7:0])}):((control_194_10)?({(operation_194_1699[7:0])}):((control_194_19)?({(operation_194_2142[7:0])}):((control_194_28)?({(operation_194_2571[7:0])}):((control_194_21)?({(operation_194_2990[7:0])}):((control_194_37)?({(operation_194_3004[7:0])}):((control_194_46)?({(operation_194_3429[7:0])}):((control_194_55)?({(operation_194_3858[7:0])}):((control_194_64)?({(operation_194_4287[7:0])}):((control_194_42)?({(operation_194_4706[7:0])}):((control_194_73)?({(operation_194_4716[7:0])}):((control_194_82)?({(operation_194_5145[7:0])}):(1'd0))))))))))))));
    assign lookup_sbox_29_enable = ((control_194_0)||((control_194_1)||((control_194_5)||((control_194_10)||((control_194_19)||((control_194_16)||((control_194_28)||((control_194_21)||((control_194_26)||((control_194_46)||((control_194_55)||((control_194_37)||((control_194_64)||((control_194_42)||((control_194_73)||((control_194_47)||((control_194_82)||(1'd0))))))))))))))))));
    assign lookup_sbox_29_0 = ((control_194_0)?({(operation_194_124[119:112])}):((control_194_1)?({(operation_194_87[7:0])}):((control_194_5)?({(operation_194_1797[7:0])}):((control_194_10)?({(operation_194_1717[7:0])}):((control_194_19)?({(operation_194_2144[7:0])}):((control_194_16)?({(operation_194_2561[7:0])}):((control_194_28)?({(operation_194_2573[7:0])}):((control_194_21)?({(operation_194_3084[7:0])}):((control_194_26)?({(operation_194_3513[7:0])}):((control_194_46)?({(operation_194_3431[7:0])}):((control_194_55)?({(operation_194_3860[7:0])}):((control_194_37)?({(operation_194_4277[7:0])}):((control_194_64)?({(operation_194_4289[7:0])}):((control_194_42)?({(operation_194_4800[7:0])}):((control_194_73)?({(operation_194_4718[7:0])}):((control_194_47)?({(operation_194_5259[7:0])}):((control_194_82)?({(operation_194_5147[7:0])}):(1'd0))))))))))))))))));
    assign lookup_sbox_30_enable = ((control_194_1)||((control_194_0)||((control_194_5)||((control_194_11)||((control_194_10)||((control_194_19)||((control_194_16)||((control_194_28)||((control_194_21)||((control_194_46)||((control_194_26)||((control_194_32)||((control_194_31)||((control_194_55)||((control_194_37)||((control_194_64)||((control_194_73)||((control_194_42)||((control_194_47)||((control_194_82)||(1'd0)))))))))))))))))))));
    assign lookup_sbox_30_0 = ((control_194_1)?({(operation_194_103[7:0])}):((control_194_0)?({(operation_194_124[111:104])}):((control_194_5)?({(operation_194_1825[7:0])}):((control_194_11)?({(operation_194_2132[7:0])}):((control_194_10)?({(operation_194_2226[7:0])}):((control_194_19)?({(operation_194_2128[7:0])}):((control_194_16)?({(operation_194_2655[7:0])}):((control_194_28)?({(operation_194_2557[7:0])}):((control_194_21)?({(operation_194_3112[7:0])}):((control_194_46)?({(operation_194_3415[7:0])}):((control_194_26)?({(operation_194_3541[7:0])}):((control_194_32)?({(operation_194_3848[7:0])}):((control_194_31)?({(operation_194_3942[7:0])}):((control_194_55)?({(operation_194_3844[7:0])}):((control_194_37)?({(operation_194_4371[7:0])}):((control_194_64)?({(operation_194_4273[7:0])}):((control_194_73)?({(operation_194_4702[7:0])}):((control_194_42)?({(operation_194_4828[7:0])}):((control_194_47)?({(operation_194_5257[7:0])}):((control_194_82)?({(operation_194_5131[7:0])}):(1'd0)))))))))))))))))))));
    assign lookup_sbox_31_enable = ((control_194_1)||((control_194_0)||((control_194_6)||((control_194_5)||((control_194_19)||((control_194_10)||((control_194_11)||((control_194_28)||((control_194_15)||((control_194_16)||((control_194_21)||((control_194_27)||((control_194_46)||((control_194_26)||((control_194_55)||((control_194_31)||((control_194_32)||((control_194_64)||((control_194_36)||((control_194_37)||((control_194_73)||((control_194_42)||((control_194_48)||((control_194_47)||((control_194_82)||(1'd0))))))))))))))))))))))))));
    assign lookup_sbox_31_0 = ((control_194_1)?({(operation_194_119[7:0])}):((control_194_0)?({(operation_194_124[127:120])}):((control_194_6)?({(operation_194_1703[7:0])}):((control_194_5)?({(operation_194_1827[7:0])}):((control_194_19)?({(operation_194_2146[7:0])}):((control_194_10)?({(operation_194_2254[7:0])}):((control_194_11)?({(operation_194_2256[7:0])}):((control_194_28)?({(operation_194_2575[7:0])}):((control_194_15)?({(operation_194_2683[7:0])}):((control_194_16)?({(operation_194_2685[7:0])}):((control_194_21)?({(operation_194_3114[7:0])}):((control_194_27)?({(operation_194_3419[7:0])}):((control_194_46)?({(operation_194_3433[7:0])}):((control_194_26)?({(operation_194_3543[7:0])}):((control_194_55)?({(operation_194_3862[7:0])}):((control_194_31)?({(operation_194_3970[7:0])}):((control_194_32)?({(operation_194_3972[7:0])}):((control_194_64)?({(operation_194_4291[7:0])}):((control_194_36)?({(operation_194_4399[7:0])}):((control_194_37)?({(operation_194_4401[7:0])}):((control_194_73)?({(operation_194_4720[7:0])}):((control_194_42)?({(operation_194_4830[7:0])}):((control_194_48)?({(operation_194_5135[7:0])}):((control_194_47)?({(operation_194_5229[7:0])}):((control_194_82)?({(operation_194_5149[7:0])}):(1'd0))))))))))))))))))))))))));
    assign input_key_194 = ((start)?(key):(input_key_194_follow));
    assign input_in_194 = ((start)?(in):(input_in_194_follow));
    assign return_194 = ({(operation_194_1569[7:0]),(operation_194_1577[7:0]),(operation_194_1585[7:0]),(operation_194_1593[7:0]),(operation_194_1601[7:0]),(operation_194_1609[7:0]),(operation_194_1617[7:0]),(operation_194_1625[7:0]),(operation_194_1633[7:0]),(operation_194_1641[7:0]),(operation_194_1649[7:0]),(operation_194_1657[7:0]),(operation_194_1665[7:0]),(operation_194_1673[7:0]),(operation_194_1681[7:0]),(operation_194_1689[7:0])});
    assign operation_194_1665 = (operation_194_1664);
    assign operation_194_1663 = ({(operation_194_1537[7:0])});
    assign operation_194_1537 = (operation_194_1536);
    assign operation_194_1633 = (operation_194_1632);
    assign operation_194_1681 = (operation_194_1680);
    assign operation_194_1679 = ({(operation_194_1553[7:0])});
    assign operation_194_1535 = ({(operation_194_1505[7:0])});
    assign operation_194_1673 = (operation_194_1672);
    assign operation_194_1689 = (operation_194_1688);
    assign operation_194_1687 = ({(operation_194_1561[7:0])});
    assign operation_194_1671 = ({(operation_194_1545[7:0])});
    assign operation_194_1505 = (operation_194_1504);
    assign operation_194_1553 = (operation_194_1552);
    assign operation_194_1601 = (operation_194_1600);
    assign operation_194_1649 = (operation_194_1648);
    assign operation_194_1551 = ({(operation_194_1521[7:0])});
    assign operation_194_1503 = ({(operation_194_1473[7:0])});
    assign operation_194_1545 = (operation_194_1544);
    assign operation_194_1561 = (operation_194_1560);
    assign operation_194_1641 = (operation_194_1640);
    assign operation_194_1657 = (operation_194_1656);
    assign operation_194_1559 = ({(operation_194_1529[7:0])});
    assign operation_194_1543 = ({(operation_194_1513[7:0])});
    assign operation_194_1473 = (operation_194_1472);
    assign operation_194_1521 = (operation_194_1520);
    assign operation_194_1569 = (operation_194_1568);
    assign operation_194_1617 = (operation_194_1616);
    assign operation_194_1519 = ({(operation_194_1489[7:0])});
    assign operation_194_1471 = ({(operation_194_1441[7:0])});
    assign operation_194_1513 = (operation_194_1512);
    assign operation_194_1529 = (operation_194_1528);
    assign operation_194_1609 = (operation_194_1608);
    assign operation_194_1625 = (operation_194_1624);
    assign operation_194_1527 = ({(operation_194_1497[7:0])});
    assign operation_194_1511 = ({(operation_194_1481[7:0])});
    assign operation_194_1441 = (operation_194_1440);
    assign operation_194_1489 = (operation_194_1488);
    assign operation_194_1585 = (operation_194_1584);
    assign operation_194_1487 = ({(operation_194_1457[7:0])});
    assign operation_194_1439 = ({(operation_194_1433[7:0])});
    assign operation_194_1433 = (operation_194_1432);
    assign operation_194_1481 = (operation_194_1480);
    assign operation_194_1497 = (operation_194_1496);
    assign operation_194_1577 = (operation_194_1576);
    assign operation_194_1593 = (operation_194_1592);
    assign operation_194_1495 = ({(operation_194_1465[7:0])});
    assign operation_194_1479 = ({(operation_194_1449[7:0])});
    assign operation_194_1428 = ({(operation_194_1408[7:0])});
    assign operation_194_1457 = (operation_194_1456);
    assign operation_194_1455 = ({(operation_194_1418[7:0])});
    assign operation_194_1449 = (operation_194_1448);
    assign operation_194_1465 = (operation_194_1464);
    assign operation_194_1685 = ({(operation_194_1323[7:0])});
    assign operation_194_1669 = ({(operation_194_1273[7:0])});
    assign operation_194_1653 = ({(operation_194_1303[7:0])});
    assign operation_194_1637 = ({(operation_194_1333[7:0])});
    assign operation_194_1621 = ({(operation_194_1283[7:0])});
    assign operation_194_1605 = ({(operation_194_1313[7:0])});
    assign operation_194_1589 = ({(operation_194_1343[7:0])});
    assign operation_194_1573 = ({(operation_194_1293[7:0])});
    assign operation_194_1463 = ({(operation_194_1423[7:0])});
    assign operation_194_1447 = ({(operation_194_1413[7:0])});
    assign operation_194_1677 = ({(operation_194_1298[7:0])});
    assign operation_194_1661 = ({(operation_194_1328[7:0])});
    assign operation_194_1645 = ({(operation_194_1278[7:0])});
    assign operation_194_1629 = ({(operation_194_1308[7:0])});
    assign operation_194_1613 = ({(operation_194_1338[7:0])});
    assign operation_194_1597 = ({(operation_194_1288[7:0])});
    assign operation_194_1581 = ({(operation_194_1318[7:0])});
    assign operation_194_1565 = ({(operation_194_1268[7:0])});
    assign operation_194_1338 = ((control_194_83)?(lookup_sbox_31_output):(operation_194_1338_latch));
    assign operation_194_1328 = ((control_194_83)?(lookup_sbox_30_output):(operation_194_1328_latch));
    assign operation_194_1318 = ((control_194_83)?(lookup_sbox_29_output):(operation_194_1318_latch));
    assign operation_194_1308 = ((control_194_83)?(lookup_sbox_28_output):(operation_194_1308_latch));
    assign operation_194_1298 = ((control_194_83)?(lookup_sbox_27_output):(operation_194_1298_latch));
    assign operation_194_1288 = ((control_194_83)?(lookup_sbox_26_output):(operation_194_1288_latch));
    assign operation_194_1278 = ((control_194_83)?(lookup_sbox_25_output):(operation_194_1278_latch));
    assign operation_194_1268 = ((control_194_83)?(lookup_sbox_24_output):(operation_194_1268_latch));
    assign operation_194_1273 = ((control_194_83)?(lookup_sbox_23_output):(operation_194_1273_latch));
    assign operation_194_1283 = ((control_194_83)?(lookup_sbox_22_output):(operation_194_1283_latch));
    assign operation_194_1293 = ((control_194_83)?(lookup_sbox_21_output):(operation_194_1293_latch));
    assign operation_194_1303 = ((control_194_83)?(lookup_sbox_20_output):(operation_194_1303_latch));
    assign operation_194_1313 = ((control_194_83)?(lookup_sbox_19_output):(operation_194_1313_latch));
    assign operation_194_1323 = ((control_194_83)?(lookup_sbox_18_output):(operation_194_1323_latch));
    assign operation_194_1333 = ((control_194_83)?(lookup_sbox_17_output):(operation_194_1333_latch));
    assign operation_194_1343 = ((control_194_83)?(lookup_sbox_16_output):(operation_194_1343_latch));
    assign operation_194_1413 = ((control_194_48)?(lookup_sbox_31_output):(operation_194_1413_latch));
    assign operation_194_1423 = ((control_194_49)?(lookup_sbox_31_output):(operation_194_1423_latch));
    assign operation_194_1408 = ((control_194_48)?(lookup_sbox_30_output):(operation_194_1408_latch));
    assign operation_194_1418 = ((control_194_48)?(lookup_sbox_29_output):(operation_194_1418_latch));
    assign operation_194_5131 = (operation_194_5132);
    assign operation_194_5133 = ({(operation_194_5135[7:0])});
    assign operation_194_5135 = (operation_194_5136);
    assign operation_194_5137 = (operation_194_5138);
    assign operation_194_5139 = (operation_194_5140);
    assign operation_194_5141 = (operation_194_5142);
    assign operation_194_5143 = (operation_194_5144);
    assign operation_194_5145 = (operation_194_5146);
    assign operation_194_5147 = (operation_194_5148);
    assign operation_194_5149 = (operation_194_5150);
    assign operation_194_5151 = ({(operation_194_5229[7:0])});
    assign operation_194_5152 = ({(operation_194_5175[7:0])});
    assign operation_194_5153 = ({(operation_194_5173[7:0])});
    assign operation_194_5154 = ({(operation_194_5171[7:0])});
    assign operation_194_5155 = ({(operation_194_5169[7:0])});
    assign operation_194_5156 = ({(operation_194_5167[7:0])});
    assign operation_194_5157 = ({(operation_194_5165[7:0])});
    assign operation_194_5158 = ({(operation_194_5163[7:0])});
    assign operation_194_5159 = ({(operation_194_5161[7:0])});
    assign operation_194_5160 = ({(operation_194_5227[7:0])});
    assign operation_194_5161 = (operation_194_5162);
    assign operation_194_5163 = (operation_194_5164);
    assign operation_194_5165 = (operation_194_5166);
    assign operation_194_5167 = (operation_194_5168);
    assign operation_194_5169 = (operation_194_5170);
    assign operation_194_5171 = (operation_194_5172);
    assign operation_194_5173 = (operation_194_5174);
    assign operation_194_5175 = (operation_194_5176);
    assign operation_194_5177 = (operation_194_5178);
    assign operation_194_5179 = (operation_194_5180);
    assign operation_194_5181 = (operation_194_5182);
    assign operation_194_5183 = (operation_194_5184);
    assign operation_194_5185 = (operation_194_5186);
    assign operation_194_5187 = (operation_194_5188);
    assign operation_194_5189 = (operation_194_5190);
    assign operation_194_5191 = (operation_194_5192);
    assign operation_194_5193 = ({(operation_194_5259[7:0])});
    assign operation_194_5194 = ({(operation_194_5225[7:0])});
    assign operation_194_5195 = ({(operation_194_5257[7:0])});
    assign operation_194_5196 = ({(operation_194_5223[7:0])});
    assign operation_194_5197 = ({(operation_194_5221[7:0])});
    assign operation_194_5198 = ({(operation_194_5219[7:0])});
    assign operation_194_5199 = ({(operation_194_5217[7:0])});
    assign operation_194_5200 = ({(operation_194_5215[7:0])});
    assign operation_194_5201 = ({(operation_194_5213[7:0])});
    assign operation_194_5202 = ({(operation_194_5211[7:0])});
    assign operation_194_5203 = ({(operation_194_5255[7:0])});
    assign operation_194_5204 = ({(operation_194_5253[7:0])});
    assign operation_194_5205 = ({(operation_194_5251[7:0])});
    assign operation_194_5206 = ({(operation_194_5249[7:0])});
    assign operation_194_5207 = ({(operation_194_5247[7:0])});
    assign operation_194_5208 = ({(operation_194_5245[7:0])});
    assign operation_194_5209 = ({(operation_194_5243[7:0])});
    assign operation_194_5210 = ({(operation_194_5241[7:0])});
    assign operation_194_5211 = (operation_194_5212);
    assign operation_194_5213 = (operation_194_5214);
    assign operation_194_5215 = (operation_194_5216);
    assign operation_194_5217 = (operation_194_5218);
    assign operation_194_5219 = (operation_194_5220);
    assign operation_194_5221 = (operation_194_5222);
    assign operation_194_5223 = (operation_194_5224);
    assign operation_194_5225 = (operation_194_5226);
    assign operation_194_5227 = (operation_194_5228);
    assign operation_194_5229 = (operation_194_5230);
    assign operation_194_5231 = ({(operation_194_5289[7:0])});
    assign operation_194_5232 = ({(operation_194_5287[7:0])});
    assign operation_194_5233 = ({(operation_194_5285[7:0])});
    assign operation_194_5234 = ({(operation_194_5283[7:0])});
    assign operation_194_5235 = ({(operation_194_5281[7:0])});
    assign operation_194_5236 = ({(operation_194_5279[7:0])});
    assign operation_194_5237 = ({(operation_194_5277[7:0])});
    assign operation_194_5238 = ({(operation_194_5275[7:0])});
    assign operation_194_5239 = ({(operation_194_5273[7:0])});
    assign operation_194_5240 = ({(operation_194_5271[7:0])});
    assign operation_194_5241 = (operation_194_5242);
    assign operation_194_5243 = (operation_194_5244);
    assign operation_194_5245 = (operation_194_5246);
    assign operation_194_5247 = (operation_194_5248);
    assign operation_194_5249 = (operation_194_5250);
    assign operation_194_5251 = (operation_194_5252);
    assign operation_194_5253 = (operation_194_5254);
    assign operation_194_5255 = (operation_194_5256);
    assign operation_194_5257 = (operation_194_5258);
    assign operation_194_5259 = (operation_194_5260);
    assign operation_194_5261 = ({(operation_194_5327[7:0])});
    assign operation_194_5262 = ({(operation_194_5325[7:0])});
    assign operation_194_5263 = ({(operation_194_5322[7:0])});
    assign operation_194_5264 = ({(operation_194_5319[7:0])});
    assign operation_194_5265 = ({(operation_194_5316[7:0])});
    assign operation_194_5266 = ({(operation_194_5313[7:0])});
    assign operation_194_5267 = ({(operation_194_5310[7:0])});
    assign operation_194_5268 = ({(operation_194_5307[7:0])});
    assign operation_194_5269 = ({(operation_194_5304[7:0])});
    assign operation_194_5270 = ({(operation_194_5301[7:0])});
    assign operation_194_5271 = (operation_194_5272);
    assign operation_194_5273 = (operation_194_5274);
    assign operation_194_5275 = (operation_194_5276);
    assign operation_194_5277 = (operation_194_5278);
    assign operation_194_5279 = (operation_194_5280);
    assign operation_194_5281 = (operation_194_5282);
    assign operation_194_5283 = (operation_194_5284);
    assign operation_194_5285 = (operation_194_5286);
    assign operation_194_5287 = (operation_194_5288);
    assign operation_194_5289 = (operation_194_5290);
    assign operation_194_5291 = ({(operation_194_5389[7:0])});
    assign operation_194_5292 = ({(operation_194_5387[7:0])});
    assign operation_194_5293 = ({(operation_194_5384[7:0])});
    assign operation_194_5294 = ({(operation_194_5381[7:0])});
    assign operation_194_5295 = ({(operation_194_5378[7:0])});
    assign operation_194_5296 = ({(operation_194_5375[7:0])});
    assign operation_194_5297 = ({(operation_194_5372[7:0])});
    assign operation_194_5298 = ({(operation_194_5369[7:0])});
    assign operation_194_5299 = ({(operation_194_5366[7:0])});
    assign operation_194_5300 = ({(operation_194_5363[7:0])});
    assign operation_194_5301 = (operation_194_5302);
    assign operation_194_5304 = (operation_194_5305);
    assign operation_194_5307 = (operation_194_5308);
    assign operation_194_5310 = (operation_194_5311);
    assign operation_194_5313 = (operation_194_5314);
    assign operation_194_5316 = (operation_194_5317);
    assign operation_194_5319 = (operation_194_5320);
    assign operation_194_5322 = (operation_194_5323);
    assign operation_194_5325 = (operation_194_5326);
    assign operation_194_5327 = (operation_194_5328);
    assign operation_194_5329 = ({(operation_194_5447[7:0])});
    assign operation_194_5330 = ({(operation_194_5445[7:0])});
    assign operation_194_5334 = ({(operation_194_5437[7:0])});
    assign operation_194_5338 = ({(operation_194_5436[7:0])});
    assign operation_194_5342 = ({(operation_194_5434[7:0])});
    assign operation_194_5346 = ({(operation_194_5433[7:0])});
    assign operation_194_5350 = ({(operation_194_5431[7:0])});
    assign operation_194_5354 = ({(operation_194_5430[7:0])});
    assign operation_194_5358 = ({(operation_194_5428[7:0])});
    assign operation_194_5362 = ({(operation_194_5427[7:0])});
    assign operation_194_5363 = (operation_194_5364);
    assign operation_194_5366 = (operation_194_5367);
    assign operation_194_5369 = (operation_194_5370);
    assign operation_194_5372 = (operation_194_5373);
    assign operation_194_5375 = (operation_194_5376);
    assign operation_194_5378 = (operation_194_5379);
    assign operation_194_5381 = (operation_194_5382);
    assign operation_194_5384 = (operation_194_5385);
    assign operation_194_5387 = (operation_194_5388);
    assign operation_194_5389 = (operation_194_5390);
    assign operation_194_5391 = ({(operation_194_5478[7:0])});
    assign operation_194_5392 = ({(operation_194_5443[7:0])});
    assign operation_194_5393 = ({(operation_194_5441[7:0])});
    assign operation_194_5394 = ({(operation_194_5439[7:0])});
    assign operation_194_5398 = ({(operation_194_5472[7:0])});
    assign operation_194_5402 = ({(operation_194_5470[7:0])});
    assign operation_194_5406 = ({(operation_194_5468[7:0])});
    assign operation_194_5410 = ({(operation_194_5466[7:0])});
    assign operation_194_5414 = ({(operation_194_5464[7:0])});
    assign operation_194_5418 = ({(operation_194_5462[7:0])});
    assign operation_194_5422 = ({(operation_194_5460[7:0])});
    assign operation_194_5426 = ({(operation_194_5458[7:0])});
    assign operation_194_5427 = (operation_194_5457);
    assign operation_194_5428 = (operation_194_5429);
    assign operation_194_5430 = (operation_194_5492);
    assign operation_194_5431 = (operation_194_5432);
    assign operation_194_5433 = (operation_194_5455);
    assign operation_194_5434 = (operation_194_5435);
    assign operation_194_5436 = (operation_194_5490);
    assign operation_194_5437 = (operation_194_5438);
    assign operation_194_5439 = (operation_194_5440);
    assign operation_194_5441 = (operation_194_5442);
    assign operation_194_5443 = (operation_194_5444);
    assign operation_194_5445 = (operation_194_5446);
    assign operation_194_5447 = (operation_194_5448);
    assign operation_194_5449 = ({(operation_194_5505[7:0])});
    assign operation_194_5450 = ({(operation_194_5503[7:0])});
    assign operation_194_5451 = ({(operation_194_5522[7:0])});
    assign operation_194_5452 = ({(operation_194_5476[7:0])});
    assign operation_194_5453 = ({(operation_194_5474[7:0])});
    assign operation_194_5458 = (operation_194_5459);
    assign operation_194_5460 = (operation_194_5461);
    assign operation_194_5462 = (operation_194_5463);
    assign operation_194_5464 = (operation_194_5465);
    assign operation_194_5466 = (operation_194_5467);
    assign operation_194_5468 = (operation_194_5469);
    assign operation_194_5470 = (operation_194_5471);
    assign operation_194_5472 = (operation_194_5473);
    assign operation_194_5474 = (operation_194_5475);
    assign operation_194_5476 = (operation_194_5477);
    assign operation_194_5478 = (operation_194_5479);
    assign operation_194_5486 = ({(operation_194_5521[7:0])});
    assign operation_194_5493 = ({(operation_194_5532[7:0])});
    assign operation_194_5494 = ({(operation_194_5535[7:0])});
    assign operation_194_5495 = ({(operation_194_5534[7:0])});
    assign operation_194_5496 = ({(operation_194_5537[7:0])});
    assign operation_194_5497 = ({(operation_194_5536[7:0])});
    assign operation_194_5498 = ({(operation_194_5531[7:0])});
    assign operation_194_5499 = ({(operation_194_5538[7:0])});
    assign operation_194_5500 = ({(operation_194_5533[7:0])});
    assign operation_194_5503 = (operation_194_5504);
    assign operation_194_5505 = (operation_194_5506);
    assign operation_194_5517 = ({(operation_194_5548[7:0])});
    assign operation_194_5519 = ({(operation_194_5547[7:0])});
    assign operation_194_5521 = ((control_194_43)?(lookup_sbox_31_output):(operation_194_5521_latch));
    assign operation_194_5522 = ((control_194_43)?(lookup_sbox_30_output):(operation_194_5522_latch));
    assign operation_194_5523 = ({(operation_194_5544[7:0])});
    assign operation_194_5524 = ({(operation_194_5539[7:0])});
    assign operation_194_5525 = ({(operation_194_5542[7:0])});
    assign operation_194_5526 = ({(operation_194_5545[7:0])});
    assign operation_194_5527 = ({(operation_194_5540[7:0])});
    assign operation_194_5528 = ({(operation_194_5543[7:0])});
    assign operation_194_5529 = ({(operation_194_5546[7:0])});
    assign operation_194_5530 = ({(operation_194_5541[7:0])});
    assign operation_194_5531 = ((control_194_74)?(lookup_sbox_31_output):(operation_194_5531_latch));
    assign operation_194_5532 = ((control_194_74)?(lookup_sbox_30_output):(operation_194_5532_latch));
    assign operation_194_5533 = ((control_194_74)?(lookup_sbox_29_output):(operation_194_5533_latch));
    assign operation_194_5534 = ((control_194_74)?(lookup_sbox_28_output):(operation_194_5534_latch));
    assign operation_194_5535 = ((control_194_74)?(lookup_sbox_27_output):(operation_194_5535_latch));
    assign operation_194_5536 = ((control_194_74)?(lookup_sbox_26_output):(operation_194_5536_latch));
    assign operation_194_5537 = ((control_194_74)?(lookup_sbox_25_output):(operation_194_5537_latch));
    assign operation_194_5538 = ((control_194_74)?(lookup_sbox_24_output):(operation_194_5538_latch));
    assign operation_194_5539 = ((control_194_74)?(lookup_sbox_23_output):(operation_194_5539_latch));
    assign operation_194_5540 = ((control_194_74)?(lookup_sbox_22_output):(operation_194_5540_latch));
    assign operation_194_5541 = ((control_194_74)?(lookup_sbox_21_output):(operation_194_5541_latch));
    assign operation_194_5542 = ((control_194_74)?(lookup_sbox_20_output):(operation_194_5542_latch));
    assign operation_194_5543 = ((control_194_74)?(lookup_sbox_19_output):(operation_194_5543_latch));
    assign operation_194_5544 = ((control_194_74)?(lookup_sbox_18_output):(operation_194_5544_latch));
    assign operation_194_5545 = ((control_194_74)?(lookup_sbox_17_output):(operation_194_5545_latch));
    assign operation_194_5546 = ((control_194_74)?(lookup_sbox_16_output):(operation_194_5546_latch));
    assign operation_194_5547 = ((control_194_43)?(lookup_sbox_29_output):(operation_194_5547_latch));
    assign operation_194_5548 = ((control_194_43)?(lookup_sbox_28_output):(operation_194_5548_latch));
    assign operation_194_4702 = (operation_194_4703);
    assign operation_194_4704 = ({(operation_194_4706[7:0])});
    assign operation_194_4706 = (operation_194_4707);
    assign operation_194_4708 = (operation_194_4709);
    assign operation_194_4710 = (operation_194_4711);
    assign operation_194_4712 = (operation_194_4713);
    assign operation_194_4714 = (operation_194_4715);
    assign operation_194_4716 = (operation_194_4717);
    assign operation_194_4718 = (operation_194_4719);
    assign operation_194_4720 = (operation_194_4721);
    assign operation_194_4722 = ({(operation_194_4800[7:0])});
    assign operation_194_4723 = ({(operation_194_4746[7:0])});
    assign operation_194_4724 = ({(operation_194_4744[7:0])});
    assign operation_194_4725 = ({(operation_194_4742[7:0])});
    assign operation_194_4726 = ({(operation_194_4740[7:0])});
    assign operation_194_4727 = ({(operation_194_4738[7:0])});
    assign operation_194_4728 = ({(operation_194_4736[7:0])});
    assign operation_194_4729 = ({(operation_194_4734[7:0])});
    assign operation_194_4730 = ({(operation_194_4732[7:0])});
    assign operation_194_4731 = ({(operation_194_4798[7:0])});
    assign operation_194_4732 = (operation_194_4733);
    assign operation_194_4734 = (operation_194_4735);
    assign operation_194_4736 = (operation_194_4737);
    assign operation_194_4738 = (operation_194_4739);
    assign operation_194_4740 = (operation_194_4741);
    assign operation_194_4742 = (operation_194_4743);
    assign operation_194_4744 = (operation_194_4745);
    assign operation_194_4746 = (operation_194_4747);
    assign operation_194_4748 = (operation_194_4749);
    assign operation_194_4750 = (operation_194_4751);
    assign operation_194_4752 = (operation_194_4753);
    assign operation_194_4754 = (operation_194_4755);
    assign operation_194_4756 = (operation_194_4757);
    assign operation_194_4758 = (operation_194_4759);
    assign operation_194_4760 = (operation_194_4761);
    assign operation_194_4762 = (operation_194_4763);
    assign operation_194_4764 = ({(operation_194_4830[7:0])});
    assign operation_194_4765 = ({(operation_194_4796[7:0])});
    assign operation_194_4766 = ({(operation_194_4828[7:0])});
    assign operation_194_4767 = ({(operation_194_4794[7:0])});
    assign operation_194_4768 = ({(operation_194_4792[7:0])});
    assign operation_194_4769 = ({(operation_194_4790[7:0])});
    assign operation_194_4770 = ({(operation_194_4788[7:0])});
    assign operation_194_4771 = ({(operation_194_4786[7:0])});
    assign operation_194_4772 = ({(operation_194_4784[7:0])});
    assign operation_194_4773 = ({(operation_194_4782[7:0])});
    assign operation_194_4774 = ({(operation_194_4826[7:0])});
    assign operation_194_4775 = ({(operation_194_4824[7:0])});
    assign operation_194_4776 = ({(operation_194_4822[7:0])});
    assign operation_194_4777 = ({(operation_194_4820[7:0])});
    assign operation_194_4778 = ({(operation_194_4818[7:0])});
    assign operation_194_4779 = ({(operation_194_4816[7:0])});
    assign operation_194_4780 = ({(operation_194_4814[7:0])});
    assign operation_194_4781 = ({(operation_194_4812[7:0])});
    assign operation_194_4782 = (operation_194_4783);
    assign operation_194_4784 = (operation_194_4785);
    assign operation_194_4786 = (operation_194_4787);
    assign operation_194_4788 = (operation_194_4789);
    assign operation_194_4790 = (operation_194_4791);
    assign operation_194_4792 = (operation_194_4793);
    assign operation_194_4794 = (operation_194_4795);
    assign operation_194_4796 = (operation_194_4797);
    assign operation_194_4798 = (operation_194_4799);
    assign operation_194_4800 = (operation_194_4801);
    assign operation_194_4802 = ({(operation_194_4860[7:0])});
    assign operation_194_4803 = ({(operation_194_4858[7:0])});
    assign operation_194_4804 = ({(operation_194_4856[7:0])});
    assign operation_194_4805 = ({(operation_194_4854[7:0])});
    assign operation_194_4806 = ({(operation_194_4852[7:0])});
    assign operation_194_4807 = ({(operation_194_4850[7:0])});
    assign operation_194_4808 = ({(operation_194_4848[7:0])});
    assign operation_194_4809 = ({(operation_194_4846[7:0])});
    assign operation_194_4810 = ({(operation_194_4844[7:0])});
    assign operation_194_4811 = ({(operation_194_4842[7:0])});
    assign operation_194_4812 = (operation_194_4813);
    assign operation_194_4814 = (operation_194_4815);
    assign operation_194_4816 = (operation_194_4817);
    assign operation_194_4818 = (operation_194_4819);
    assign operation_194_4820 = (operation_194_4821);
    assign operation_194_4822 = (operation_194_4823);
    assign operation_194_4824 = (operation_194_4825);
    assign operation_194_4826 = (operation_194_4827);
    assign operation_194_4828 = (operation_194_4829);
    assign operation_194_4830 = (operation_194_4831);
    assign operation_194_4832 = ({(operation_194_4898[7:0])});
    assign operation_194_4833 = ({(operation_194_4896[7:0])});
    assign operation_194_4834 = ({(operation_194_4893[7:0])});
    assign operation_194_4835 = ({(operation_194_4890[7:0])});
    assign operation_194_4836 = ({(operation_194_4887[7:0])});
    assign operation_194_4837 = ({(operation_194_4884[7:0])});
    assign operation_194_4838 = ({(operation_194_4881[7:0])});
    assign operation_194_4839 = ({(operation_194_4878[7:0])});
    assign operation_194_4840 = ({(operation_194_4875[7:0])});
    assign operation_194_4841 = ({(operation_194_4872[7:0])});
    assign operation_194_4842 = (operation_194_4843);
    assign operation_194_4844 = (operation_194_4845);
    assign operation_194_4846 = (operation_194_4847);
    assign operation_194_4848 = (operation_194_4849);
    assign operation_194_4850 = (operation_194_4851);
    assign operation_194_4852 = (operation_194_4853);
    assign operation_194_4854 = (operation_194_4855);
    assign operation_194_4856 = (operation_194_4857);
    assign operation_194_4858 = (operation_194_4859);
    assign operation_194_4860 = (operation_194_4861);
    assign operation_194_4862 = ({(operation_194_4960[7:0])});
    assign operation_194_4863 = ({(operation_194_4958[7:0])});
    assign operation_194_4864 = ({(operation_194_4955[7:0])});
    assign operation_194_4865 = ({(operation_194_4952[7:0])});
    assign operation_194_4866 = ({(operation_194_4949[7:0])});
    assign operation_194_4867 = ({(operation_194_4946[7:0])});
    assign operation_194_4868 = ({(operation_194_4943[7:0])});
    assign operation_194_4869 = ({(operation_194_4940[7:0])});
    assign operation_194_4870 = ({(operation_194_4937[7:0])});
    assign operation_194_4871 = ({(operation_194_4934[7:0])});
    assign operation_194_4872 = (operation_194_4873);
    assign operation_194_4875 = (operation_194_4876);
    assign operation_194_4878 = (operation_194_4879);
    assign operation_194_4881 = (operation_194_4882);
    assign operation_194_4884 = (operation_194_4885);
    assign operation_194_4887 = (operation_194_4888);
    assign operation_194_4890 = (operation_194_4891);
    assign operation_194_4893 = (operation_194_4894);
    assign operation_194_4896 = (operation_194_4897);
    assign operation_194_4898 = (operation_194_4899);
    assign operation_194_4900 = ({(operation_194_5018[7:0])});
    assign operation_194_4901 = ({(operation_194_5016[7:0])});
    assign operation_194_4905 = ({(operation_194_5008[7:0])});
    assign operation_194_4909 = ({(operation_194_5007[7:0])});
    assign operation_194_4913 = ({(operation_194_5005[7:0])});
    assign operation_194_4917 = ({(operation_194_5004[7:0])});
    assign operation_194_4921 = ({(operation_194_5002[7:0])});
    assign operation_194_4925 = ({(operation_194_5001[7:0])});
    assign operation_194_4929 = ({(operation_194_4999[7:0])});
    assign operation_194_4933 = ({(operation_194_4998[7:0])});
    assign operation_194_4934 = (operation_194_4935);
    assign operation_194_4937 = (operation_194_4938);
    assign operation_194_4940 = (operation_194_4941);
    assign operation_194_4943 = (operation_194_4944);
    assign operation_194_4946 = (operation_194_4947);
    assign operation_194_4949 = (operation_194_4950);
    assign operation_194_4952 = (operation_194_4953);
    assign operation_194_4955 = (operation_194_4956);
    assign operation_194_4958 = (operation_194_4959);
    assign operation_194_4960 = (operation_194_4961);
    assign operation_194_4962 = ({(operation_194_5049[7:0])});
    assign operation_194_4963 = ({(operation_194_5014[7:0])});
    assign operation_194_4964 = ({(operation_194_5012[7:0])});
    assign operation_194_4965 = ({(operation_194_5010[7:0])});
    assign operation_194_4969 = ({(operation_194_5043[7:0])});
    assign operation_194_4973 = ({(operation_194_5041[7:0])});
    assign operation_194_4977 = ({(operation_194_5039[7:0])});
    assign operation_194_4981 = ({(operation_194_5037[7:0])});
    assign operation_194_4985 = ({(operation_194_5035[7:0])});
    assign operation_194_4989 = ({(operation_194_5033[7:0])});
    assign operation_194_4993 = ({(operation_194_5031[7:0])});
    assign operation_194_4997 = ({(operation_194_5029[7:0])});
    assign operation_194_4998 = (operation_194_5028);
    assign operation_194_4999 = (operation_194_5000);
    assign operation_194_5001 = (operation_194_5063);
    assign operation_194_5002 = (operation_194_5003);
    assign operation_194_5004 = (operation_194_5026);
    assign operation_194_5005 = (operation_194_5006);
    assign operation_194_5007 = (operation_194_5061);
    assign operation_194_5008 = (operation_194_5009);
    assign operation_194_5010 = (operation_194_5011);
    assign operation_194_5012 = (operation_194_5013);
    assign operation_194_5014 = (operation_194_5015);
    assign operation_194_5016 = (operation_194_5017);
    assign operation_194_5018 = (operation_194_5019);
    assign operation_194_5020 = ({(operation_194_5076[7:0])});
    assign operation_194_5021 = ({(operation_194_5074[7:0])});
    assign operation_194_5022 = ({(operation_194_5093[7:0])});
    assign operation_194_5023 = ({(operation_194_5047[7:0])});
    assign operation_194_5024 = ({(operation_194_5045[7:0])});
    assign operation_194_5029 = (operation_194_5030);
    assign operation_194_5031 = (operation_194_5032);
    assign operation_194_5033 = (operation_194_5034);
    assign operation_194_5035 = (operation_194_5036);
    assign operation_194_5037 = (operation_194_5038);
    assign operation_194_5039 = (operation_194_5040);
    assign operation_194_5041 = (operation_194_5042);
    assign operation_194_5043 = (operation_194_5044);
    assign operation_194_5045 = (operation_194_5046);
    assign operation_194_5047 = (operation_194_5048);
    assign operation_194_5049 = (operation_194_5050);
    assign operation_194_5057 = ({(operation_194_5092[7:0])});
    assign operation_194_5064 = ({(operation_194_5103[7:0])});
    assign operation_194_5065 = ({(operation_194_5106[7:0])});
    assign operation_194_5066 = ({(operation_194_5105[7:0])});
    assign operation_194_5067 = ({(operation_194_5108[7:0])});
    assign operation_194_5068 = ({(operation_194_5107[7:0])});
    assign operation_194_5069 = ({(operation_194_5102[7:0])});
    assign operation_194_5070 = ({(operation_194_5109[7:0])});
    assign operation_194_5071 = ({(operation_194_5104[7:0])});
    assign operation_194_5074 = (operation_194_5075);
    assign operation_194_5076 = (operation_194_5077);
    assign operation_194_5088 = ({(operation_194_5119[7:0])});
    assign operation_194_5090 = ({(operation_194_5118[7:0])});
    assign operation_194_5092 = ((control_194_38)?(lookup_sbox_31_output):(operation_194_5092_latch));
    assign operation_194_5093 = ((control_194_37)?(lookup_sbox_31_output):(operation_194_5093_latch));
    assign operation_194_5094 = ({(operation_194_5115[7:0])});
    assign operation_194_5095 = ({(operation_194_5110[7:0])});
    assign operation_194_5096 = ({(operation_194_5113[7:0])});
    assign operation_194_5097 = ({(operation_194_5116[7:0])});
    assign operation_194_5098 = ({(operation_194_5111[7:0])});
    assign operation_194_5099 = ({(operation_194_5114[7:0])});
    assign operation_194_5100 = ({(operation_194_5117[7:0])});
    assign operation_194_5101 = ({(operation_194_5112[7:0])});
    assign operation_194_5102 = ((control_194_65)?(lookup_sbox_31_output):(operation_194_5102_latch));
    assign operation_194_5103 = ((control_194_65)?(lookup_sbox_30_output):(operation_194_5103_latch));
    assign operation_194_5104 = ((control_194_65)?(lookup_sbox_29_output):(operation_194_5104_latch));
    assign operation_194_5105 = ((control_194_65)?(lookup_sbox_28_output):(operation_194_5105_latch));
    assign operation_194_5106 = ((control_194_65)?(lookup_sbox_27_output):(operation_194_5106_latch));
    assign operation_194_5107 = ((control_194_65)?(lookup_sbox_26_output):(operation_194_5107_latch));
    assign operation_194_5108 = ((control_194_65)?(lookup_sbox_25_output):(operation_194_5108_latch));
    assign operation_194_5109 = ((control_194_65)?(lookup_sbox_24_output):(operation_194_5109_latch));
    assign operation_194_5110 = ((control_194_65)?(lookup_sbox_23_output):(operation_194_5110_latch));
    assign operation_194_5111 = ((control_194_65)?(lookup_sbox_22_output):(operation_194_5111_latch));
    assign operation_194_5112 = ((control_194_65)?(lookup_sbox_21_output):(operation_194_5112_latch));
    assign operation_194_5113 = ((control_194_65)?(lookup_sbox_20_output):(operation_194_5113_latch));
    assign operation_194_5114 = ((control_194_65)?(lookup_sbox_19_output):(operation_194_5114_latch));
    assign operation_194_5115 = ((control_194_65)?(lookup_sbox_18_output):(operation_194_5115_latch));
    assign operation_194_5116 = ((control_194_65)?(lookup_sbox_17_output):(operation_194_5116_latch));
    assign operation_194_5117 = ((control_194_65)?(lookup_sbox_16_output):(operation_194_5117_latch));
    assign operation_194_5118 = ((control_194_38)?(lookup_sbox_30_output):(operation_194_5118_latch));
    assign operation_194_5119 = ((control_194_38)?(lookup_sbox_29_output):(operation_194_5119_latch));
    assign operation_194_4273 = (operation_194_4274);
    assign operation_194_4275 = ({(operation_194_4277[7:0])});
    assign operation_194_4277 = (operation_194_4278);
    assign operation_194_4279 = (operation_194_4280);
    assign operation_194_4281 = (operation_194_4282);
    assign operation_194_4283 = (operation_194_4284);
    assign operation_194_4285 = (operation_194_4286);
    assign operation_194_4287 = (operation_194_4288);
    assign operation_194_4289 = (operation_194_4290);
    assign operation_194_4291 = (operation_194_4292);
    assign operation_194_4293 = ({(operation_194_4371[7:0])});
    assign operation_194_4294 = ({(operation_194_4317[7:0])});
    assign operation_194_4295 = ({(operation_194_4315[7:0])});
    assign operation_194_4296 = ({(operation_194_4313[7:0])});
    assign operation_194_4297 = ({(operation_194_4311[7:0])});
    assign operation_194_4298 = ({(operation_194_4309[7:0])});
    assign operation_194_4299 = ({(operation_194_4307[7:0])});
    assign operation_194_4300 = ({(operation_194_4305[7:0])});
    assign operation_194_4301 = ({(operation_194_4303[7:0])});
    assign operation_194_4302 = ({(operation_194_4369[7:0])});
    assign operation_194_4303 = (operation_194_4304);
    assign operation_194_4305 = (operation_194_4306);
    assign operation_194_4307 = (operation_194_4308);
    assign operation_194_4309 = (operation_194_4310);
    assign operation_194_4311 = (operation_194_4312);
    assign operation_194_4313 = (operation_194_4314);
    assign operation_194_4315 = (operation_194_4316);
    assign operation_194_4317 = (operation_194_4318);
    assign operation_194_4319 = (operation_194_4320);
    assign operation_194_4321 = (operation_194_4322);
    assign operation_194_4323 = (operation_194_4324);
    assign operation_194_4325 = (operation_194_4326);
    assign operation_194_4327 = (operation_194_4328);
    assign operation_194_4329 = (operation_194_4330);
    assign operation_194_4331 = (operation_194_4332);
    assign operation_194_4333 = (operation_194_4334);
    assign operation_194_4335 = ({(operation_194_4401[7:0])});
    assign operation_194_4336 = ({(operation_194_4367[7:0])});
    assign operation_194_4337 = ({(operation_194_4399[7:0])});
    assign operation_194_4338 = ({(operation_194_4365[7:0])});
    assign operation_194_4339 = ({(operation_194_4363[7:0])});
    assign operation_194_4340 = ({(operation_194_4361[7:0])});
    assign operation_194_4341 = ({(operation_194_4359[7:0])});
    assign operation_194_4342 = ({(operation_194_4357[7:0])});
    assign operation_194_4343 = ({(operation_194_4355[7:0])});
    assign operation_194_4344 = ({(operation_194_4353[7:0])});
    assign operation_194_4345 = ({(operation_194_4397[7:0])});
    assign operation_194_4346 = ({(operation_194_4395[7:0])});
    assign operation_194_4347 = ({(operation_194_4393[7:0])});
    assign operation_194_4348 = ({(operation_194_4391[7:0])});
    assign operation_194_4349 = ({(operation_194_4389[7:0])});
    assign operation_194_4350 = ({(operation_194_4387[7:0])});
    assign operation_194_4351 = ({(operation_194_4385[7:0])});
    assign operation_194_4352 = ({(operation_194_4383[7:0])});
    assign operation_194_4353 = (operation_194_4354);
    assign operation_194_4355 = (operation_194_4356);
    assign operation_194_4357 = (operation_194_4358);
    assign operation_194_4359 = (operation_194_4360);
    assign operation_194_4361 = (operation_194_4362);
    assign operation_194_4363 = (operation_194_4364);
    assign operation_194_4365 = (operation_194_4366);
    assign operation_194_4367 = (operation_194_4368);
    assign operation_194_4369 = (operation_194_4370);
    assign operation_194_4371 = (operation_194_4372);
    assign operation_194_4373 = ({(operation_194_4431[7:0])});
    assign operation_194_4374 = ({(operation_194_4429[7:0])});
    assign operation_194_4375 = ({(operation_194_4427[7:0])});
    assign operation_194_4376 = ({(operation_194_4425[7:0])});
    assign operation_194_4377 = ({(operation_194_4423[7:0])});
    assign operation_194_4378 = ({(operation_194_4421[7:0])});
    assign operation_194_4379 = ({(operation_194_4419[7:0])});
    assign operation_194_4380 = ({(operation_194_4417[7:0])});
    assign operation_194_4381 = ({(operation_194_4415[7:0])});
    assign operation_194_4382 = ({(operation_194_4413[7:0])});
    assign operation_194_4383 = (operation_194_4384);
    assign operation_194_4385 = (operation_194_4386);
    assign operation_194_4387 = (operation_194_4388);
    assign operation_194_4389 = (operation_194_4390);
    assign operation_194_4391 = (operation_194_4392);
    assign operation_194_4393 = (operation_194_4394);
    assign operation_194_4395 = (operation_194_4396);
    assign operation_194_4397 = (operation_194_4398);
    assign operation_194_4399 = (operation_194_4400);
    assign operation_194_4401 = (operation_194_4402);
    assign operation_194_4403 = ({(operation_194_4469[7:0])});
    assign operation_194_4404 = ({(operation_194_4467[7:0])});
    assign operation_194_4405 = ({(operation_194_4464[7:0])});
    assign operation_194_4406 = ({(operation_194_4461[7:0])});
    assign operation_194_4407 = ({(operation_194_4458[7:0])});
    assign operation_194_4408 = ({(operation_194_4455[7:0])});
    assign operation_194_4409 = ({(operation_194_4452[7:0])});
    assign operation_194_4410 = ({(operation_194_4449[7:0])});
    assign operation_194_4411 = ({(operation_194_4446[7:0])});
    assign operation_194_4412 = ({(operation_194_4443[7:0])});
    assign operation_194_4413 = (operation_194_4414);
    assign operation_194_4415 = (operation_194_4416);
    assign operation_194_4417 = (operation_194_4418);
    assign operation_194_4419 = (operation_194_4420);
    assign operation_194_4421 = (operation_194_4422);
    assign operation_194_4423 = (operation_194_4424);
    assign operation_194_4425 = (operation_194_4426);
    assign operation_194_4427 = (operation_194_4428);
    assign operation_194_4429 = (operation_194_4430);
    assign operation_194_4431 = (operation_194_4432);
    assign operation_194_4433 = ({(operation_194_4531[7:0])});
    assign operation_194_4434 = ({(operation_194_4529[7:0])});
    assign operation_194_4435 = ({(operation_194_4526[7:0])});
    assign operation_194_4436 = ({(operation_194_4523[7:0])});
    assign operation_194_4437 = ({(operation_194_4520[7:0])});
    assign operation_194_4438 = ({(operation_194_4517[7:0])});
    assign operation_194_4439 = ({(operation_194_4514[7:0])});
    assign operation_194_4440 = ({(operation_194_4511[7:0])});
    assign operation_194_4441 = ({(operation_194_4508[7:0])});
    assign operation_194_4442 = ({(operation_194_4505[7:0])});
    assign operation_194_4443 = (operation_194_4444);
    assign operation_194_4446 = (operation_194_4447);
    assign operation_194_4449 = (operation_194_4450);
    assign operation_194_4452 = (operation_194_4453);
    assign operation_194_4455 = (operation_194_4456);
    assign operation_194_4458 = (operation_194_4459);
    assign operation_194_4461 = (operation_194_4462);
    assign operation_194_4464 = (operation_194_4465);
    assign operation_194_4467 = (operation_194_4468);
    assign operation_194_4469 = (operation_194_4470);
    assign operation_194_4471 = ({(operation_194_4589[7:0])});
    assign operation_194_4472 = ({(operation_194_4587[7:0])});
    assign operation_194_4476 = ({(operation_194_4579[7:0])});
    assign operation_194_4480 = ({(operation_194_4578[7:0])});
    assign operation_194_4484 = ({(operation_194_4576[7:0])});
    assign operation_194_4488 = ({(operation_194_4575[7:0])});
    assign operation_194_4492 = ({(operation_194_4573[7:0])});
    assign operation_194_4496 = ({(operation_194_4572[7:0])});
    assign operation_194_4500 = ({(operation_194_4570[7:0])});
    assign operation_194_4504 = ({(operation_194_4569[7:0])});
    assign operation_194_4505 = (operation_194_4506);
    assign operation_194_4508 = (operation_194_4509);
    assign operation_194_4511 = (operation_194_4512);
    assign operation_194_4514 = (operation_194_4515);
    assign operation_194_4517 = (operation_194_4518);
    assign operation_194_4520 = (operation_194_4521);
    assign operation_194_4523 = (operation_194_4524);
    assign operation_194_4526 = (operation_194_4527);
    assign operation_194_4529 = (operation_194_4530);
    assign operation_194_4531 = (operation_194_4532);
    assign operation_194_4533 = ({(operation_194_4620[7:0])});
    assign operation_194_4534 = ({(operation_194_4585[7:0])});
    assign operation_194_4535 = ({(operation_194_4583[7:0])});
    assign operation_194_4536 = ({(operation_194_4581[7:0])});
    assign operation_194_4540 = ({(operation_194_4614[7:0])});
    assign operation_194_4544 = ({(operation_194_4612[7:0])});
    assign operation_194_4548 = ({(operation_194_4610[7:0])});
    assign operation_194_4552 = ({(operation_194_4608[7:0])});
    assign operation_194_4556 = ({(operation_194_4606[7:0])});
    assign operation_194_4560 = ({(operation_194_4604[7:0])});
    assign operation_194_4564 = ({(operation_194_4602[7:0])});
    assign operation_194_4568 = ({(operation_194_4600[7:0])});
    assign operation_194_4569 = (operation_194_4599);
    assign operation_194_4570 = (operation_194_4571);
    assign operation_194_4572 = (operation_194_4634);
    assign operation_194_4573 = (operation_194_4574);
    assign operation_194_4575 = (operation_194_4597);
    assign operation_194_4576 = (operation_194_4577);
    assign operation_194_4578 = (operation_194_4632);
    assign operation_194_4579 = (operation_194_4580);
    assign operation_194_4581 = (operation_194_4582);
    assign operation_194_4583 = (operation_194_4584);
    assign operation_194_4585 = (operation_194_4586);
    assign operation_194_4587 = (operation_194_4588);
    assign operation_194_4589 = (operation_194_4590);
    assign operation_194_4591 = ({(operation_194_4647[7:0])});
    assign operation_194_4592 = ({(operation_194_4645[7:0])});
    assign operation_194_4593 = ({(operation_194_4664[7:0])});
    assign operation_194_4594 = ({(operation_194_4618[7:0])});
    assign operation_194_4595 = ({(operation_194_4616[7:0])});
    assign operation_194_4600 = (operation_194_4601);
    assign operation_194_4602 = (operation_194_4603);
    assign operation_194_4604 = (operation_194_4605);
    assign operation_194_4606 = (operation_194_4607);
    assign operation_194_4608 = (operation_194_4609);
    assign operation_194_4610 = (operation_194_4611);
    assign operation_194_4612 = (operation_194_4613);
    assign operation_194_4614 = (operation_194_4615);
    assign operation_194_4616 = (operation_194_4617);
    assign operation_194_4618 = (operation_194_4619);
    assign operation_194_4620 = (operation_194_4621);
    assign operation_194_4628 = ({(operation_194_4663[7:0])});
    assign operation_194_4635 = ({(operation_194_4674[7:0])});
    assign operation_194_4636 = ({(operation_194_4677[7:0])});
    assign operation_194_4637 = ({(operation_194_4676[7:0])});
    assign operation_194_4638 = ({(operation_194_4679[7:0])});
    assign operation_194_4639 = ({(operation_194_4678[7:0])});
    assign operation_194_4640 = ({(operation_194_4673[7:0])});
    assign operation_194_4641 = ({(operation_194_4680[7:0])});
    assign operation_194_4642 = ({(operation_194_4675[7:0])});
    assign operation_194_4645 = (operation_194_4646);
    assign operation_194_4647 = (operation_194_4648);
    assign operation_194_4659 = ({(operation_194_4690[7:0])});
    assign operation_194_4661 = ({(operation_194_4689[7:0])});
    assign operation_194_4663 = ((control_194_33)?(lookup_sbox_31_output):(operation_194_4663_latch));
    assign operation_194_4664 = ((control_194_32)?(lookup_sbox_31_output):(operation_194_4664_latch));
    assign operation_194_4665 = ({(operation_194_4686[7:0])});
    assign operation_194_4666 = ({(operation_194_4681[7:0])});
    assign operation_194_4667 = ({(operation_194_4684[7:0])});
    assign operation_194_4668 = ({(operation_194_4687[7:0])});
    assign operation_194_4669 = ({(operation_194_4682[7:0])});
    assign operation_194_4670 = ({(operation_194_4685[7:0])});
    assign operation_194_4671 = ({(operation_194_4688[7:0])});
    assign operation_194_4672 = ({(operation_194_4683[7:0])});
    assign operation_194_4673 = ((control_194_56)?(lookup_sbox_31_output):(operation_194_4673_latch));
    assign operation_194_4674 = ((control_194_56)?(lookup_sbox_30_output):(operation_194_4674_latch));
    assign operation_194_4675 = ((control_194_56)?(lookup_sbox_29_output):(operation_194_4675_latch));
    assign operation_194_4676 = ((control_194_56)?(lookup_sbox_28_output):(operation_194_4676_latch));
    assign operation_194_4677 = ((control_194_56)?(lookup_sbox_27_output):(operation_194_4677_latch));
    assign operation_194_4678 = ((control_194_56)?(lookup_sbox_26_output):(operation_194_4678_latch));
    assign operation_194_4679 = ((control_194_56)?(lookup_sbox_25_output):(operation_194_4679_latch));
    assign operation_194_4680 = ((control_194_56)?(lookup_sbox_24_output):(operation_194_4680_latch));
    assign operation_194_4681 = ((control_194_56)?(lookup_sbox_23_output):(operation_194_4681_latch));
    assign operation_194_4682 = ((control_194_56)?(lookup_sbox_22_output):(operation_194_4682_latch));
    assign operation_194_4683 = ((control_194_56)?(lookup_sbox_21_output):(operation_194_4683_latch));
    assign operation_194_4684 = ((control_194_56)?(lookup_sbox_20_output):(operation_194_4684_latch));
    assign operation_194_4685 = ((control_194_56)?(lookup_sbox_19_output):(operation_194_4685_latch));
    assign operation_194_4686 = ((control_194_56)?(lookup_sbox_18_output):(operation_194_4686_latch));
    assign operation_194_4687 = ((control_194_56)?(lookup_sbox_17_output):(operation_194_4687_latch));
    assign operation_194_4688 = ((control_194_56)?(lookup_sbox_16_output):(operation_194_4688_latch));
    assign operation_194_4689 = ((control_194_32)?(lookup_sbox_30_output):(operation_194_4689_latch));
    assign operation_194_4690 = ((control_194_33)?(lookup_sbox_30_output):(operation_194_4690_latch));
    assign operation_194_3844 = (operation_194_3845);
    assign operation_194_3846 = ({(operation_194_3848[7:0])});
    assign operation_194_3848 = (operation_194_3849);
    assign operation_194_3850 = (operation_194_3851);
    assign operation_194_3852 = (operation_194_3853);
    assign operation_194_3854 = (operation_194_3855);
    assign operation_194_3856 = (operation_194_3857);
    assign operation_194_3858 = (operation_194_3859);
    assign operation_194_3860 = (operation_194_3861);
    assign operation_194_3862 = (operation_194_3863);
    assign operation_194_3864 = ({(operation_194_3942[7:0])});
    assign operation_194_3865 = ({(operation_194_3888[7:0])});
    assign operation_194_3866 = ({(operation_194_3886[7:0])});
    assign operation_194_3867 = ({(operation_194_3884[7:0])});
    assign operation_194_3868 = ({(operation_194_3882[7:0])});
    assign operation_194_3869 = ({(operation_194_3880[7:0])});
    assign operation_194_3870 = ({(operation_194_3878[7:0])});
    assign operation_194_3871 = ({(operation_194_3876[7:0])});
    assign operation_194_3872 = ({(operation_194_3874[7:0])});
    assign operation_194_3873 = ({(operation_194_3940[7:0])});
    assign operation_194_3874 = (operation_194_3875);
    assign operation_194_3876 = (operation_194_3877);
    assign operation_194_3878 = (operation_194_3879);
    assign operation_194_3880 = (operation_194_3881);
    assign operation_194_3882 = (operation_194_3883);
    assign operation_194_3884 = (operation_194_3885);
    assign operation_194_3886 = (operation_194_3887);
    assign operation_194_3888 = (operation_194_3889);
    assign operation_194_3890 = (operation_194_3891);
    assign operation_194_3892 = (operation_194_3893);
    assign operation_194_3894 = (operation_194_3895);
    assign operation_194_3896 = (operation_194_3897);
    assign operation_194_3898 = (operation_194_3899);
    assign operation_194_3900 = (operation_194_3901);
    assign operation_194_3902 = (operation_194_3903);
    assign operation_194_3904 = (operation_194_3905);
    assign operation_194_3906 = ({(operation_194_3972[7:0])});
    assign operation_194_3907 = ({(operation_194_3938[7:0])});
    assign operation_194_3908 = ({(operation_194_3970[7:0])});
    assign operation_194_3909 = ({(operation_194_3936[7:0])});
    assign operation_194_3910 = ({(operation_194_3934[7:0])});
    assign operation_194_3911 = ({(operation_194_3932[7:0])});
    assign operation_194_3912 = ({(operation_194_3930[7:0])});
    assign operation_194_3913 = ({(operation_194_3928[7:0])});
    assign operation_194_3914 = ({(operation_194_3926[7:0])});
    assign operation_194_3915 = ({(operation_194_3924[7:0])});
    assign operation_194_3916 = ({(operation_194_3968[7:0])});
    assign operation_194_3917 = ({(operation_194_3966[7:0])});
    assign operation_194_3918 = ({(operation_194_3964[7:0])});
    assign operation_194_3919 = ({(operation_194_3962[7:0])});
    assign operation_194_3920 = ({(operation_194_3960[7:0])});
    assign operation_194_3921 = ({(operation_194_3958[7:0])});
    assign operation_194_3922 = ({(operation_194_3956[7:0])});
    assign operation_194_3923 = ({(operation_194_3954[7:0])});
    assign operation_194_3924 = (operation_194_3925);
    assign operation_194_3926 = (operation_194_3927);
    assign operation_194_3928 = (operation_194_3929);
    assign operation_194_3930 = (operation_194_3931);
    assign operation_194_3932 = (operation_194_3933);
    assign operation_194_3934 = (operation_194_3935);
    assign operation_194_3936 = (operation_194_3937);
    assign operation_194_3938 = (operation_194_3939);
    assign operation_194_3940 = (operation_194_3941);
    assign operation_194_3942 = (operation_194_3943);
    assign operation_194_3944 = ({(operation_194_4002[7:0])});
    assign operation_194_3945 = ({(operation_194_4000[7:0])});
    assign operation_194_3946 = ({(operation_194_3998[7:0])});
    assign operation_194_3947 = ({(operation_194_3996[7:0])});
    assign operation_194_3948 = ({(operation_194_3994[7:0])});
    assign operation_194_3949 = ({(operation_194_3992[7:0])});
    assign operation_194_3950 = ({(operation_194_3990[7:0])});
    assign operation_194_3951 = ({(operation_194_3988[7:0])});
    assign operation_194_3952 = ({(operation_194_3986[7:0])});
    assign operation_194_3953 = ({(operation_194_3984[7:0])});
    assign operation_194_3954 = (operation_194_3955);
    assign operation_194_3956 = (operation_194_3957);
    assign operation_194_3958 = (operation_194_3959);
    assign operation_194_3960 = (operation_194_3961);
    assign operation_194_3962 = (operation_194_3963);
    assign operation_194_3964 = (operation_194_3965);
    assign operation_194_3966 = (operation_194_3967);
    assign operation_194_3968 = (operation_194_3969);
    assign operation_194_3970 = (operation_194_3971);
    assign operation_194_3972 = (operation_194_3973);
    assign operation_194_3974 = ({(operation_194_4040[7:0])});
    assign operation_194_3975 = ({(operation_194_4038[7:0])});
    assign operation_194_3976 = ({(operation_194_4035[7:0])});
    assign operation_194_3977 = ({(operation_194_4032[7:0])});
    assign operation_194_3978 = ({(operation_194_4029[7:0])});
    assign operation_194_3979 = ({(operation_194_4026[7:0])});
    assign operation_194_3980 = ({(operation_194_4023[7:0])});
    assign operation_194_3981 = ({(operation_194_4020[7:0])});
    assign operation_194_3982 = ({(operation_194_4017[7:0])});
    assign operation_194_3983 = ({(operation_194_4014[7:0])});
    assign operation_194_3984 = (operation_194_3985);
    assign operation_194_3986 = (operation_194_3987);
    assign operation_194_3988 = (operation_194_3989);
    assign operation_194_3990 = (operation_194_3991);
    assign operation_194_3992 = (operation_194_3993);
    assign operation_194_3994 = (operation_194_3995);
    assign operation_194_3996 = (operation_194_3997);
    assign operation_194_3998 = (operation_194_3999);
    assign operation_194_4000 = (operation_194_4001);
    assign operation_194_4002 = (operation_194_4003);
    assign operation_194_4004 = ({(operation_194_4102[7:0])});
    assign operation_194_4005 = ({(operation_194_4100[7:0])});
    assign operation_194_4006 = ({(operation_194_4097[7:0])});
    assign operation_194_4007 = ({(operation_194_4094[7:0])});
    assign operation_194_4008 = ({(operation_194_4091[7:0])});
    assign operation_194_4009 = ({(operation_194_4088[7:0])});
    assign operation_194_4010 = ({(operation_194_4085[7:0])});
    assign operation_194_4011 = ({(operation_194_4082[7:0])});
    assign operation_194_4012 = ({(operation_194_4079[7:0])});
    assign operation_194_4013 = ({(operation_194_4076[7:0])});
    assign operation_194_4014 = (operation_194_4015);
    assign operation_194_4017 = (operation_194_4018);
    assign operation_194_4020 = (operation_194_4021);
    assign operation_194_4023 = (operation_194_4024);
    assign operation_194_4026 = (operation_194_4027);
    assign operation_194_4029 = (operation_194_4030);
    assign operation_194_4032 = (operation_194_4033);
    assign operation_194_4035 = (operation_194_4036);
    assign operation_194_4038 = (operation_194_4039);
    assign operation_194_4040 = (operation_194_4041);
    assign operation_194_4042 = ({(operation_194_4160[7:0])});
    assign operation_194_4043 = ({(operation_194_4158[7:0])});
    assign operation_194_4047 = ({(operation_194_4150[7:0])});
    assign operation_194_4051 = ({(operation_194_4149[7:0])});
    assign operation_194_4055 = ({(operation_194_4147[7:0])});
    assign operation_194_4059 = ({(operation_194_4146[7:0])});
    assign operation_194_4063 = ({(operation_194_4144[7:0])});
    assign operation_194_4067 = ({(operation_194_4143[7:0])});
    assign operation_194_4071 = ({(operation_194_4141[7:0])});
    assign operation_194_4075 = ({(operation_194_4140[7:0])});
    assign operation_194_4076 = (operation_194_4077);
    assign operation_194_4079 = (operation_194_4080);
    assign operation_194_4082 = (operation_194_4083);
    assign operation_194_4085 = (operation_194_4086);
    assign operation_194_4088 = (operation_194_4089);
    assign operation_194_4091 = (operation_194_4092);
    assign operation_194_4094 = (operation_194_4095);
    assign operation_194_4097 = (operation_194_4098);
    assign operation_194_4100 = (operation_194_4101);
    assign operation_194_4102 = (operation_194_4103);
    assign operation_194_4104 = ({(operation_194_4191[7:0])});
    assign operation_194_4105 = ({(operation_194_4156[7:0])});
    assign operation_194_4106 = ({(operation_194_4154[7:0])});
    assign operation_194_4107 = ({(operation_194_4152[7:0])});
    assign operation_194_4111 = ({(operation_194_4185[7:0])});
    assign operation_194_4115 = ({(operation_194_4183[7:0])});
    assign operation_194_4119 = ({(operation_194_4181[7:0])});
    assign operation_194_4123 = ({(operation_194_4179[7:0])});
    assign operation_194_4127 = ({(operation_194_4177[7:0])});
    assign operation_194_4131 = ({(operation_194_4175[7:0])});
    assign operation_194_4135 = ({(operation_194_4173[7:0])});
    assign operation_194_4139 = ({(operation_194_4171[7:0])});
    assign operation_194_4140 = (operation_194_4170);
    assign operation_194_4141 = (operation_194_4142);
    assign operation_194_4143 = (operation_194_4205);
    assign operation_194_4144 = (operation_194_4145);
    assign operation_194_4146 = (operation_194_4168);
    assign operation_194_4147 = (operation_194_4148);
    assign operation_194_4149 = (operation_194_4203);
    assign operation_194_4150 = (operation_194_4151);
    assign operation_194_4152 = (operation_194_4153);
    assign operation_194_4154 = (operation_194_4155);
    assign operation_194_4156 = (operation_194_4157);
    assign operation_194_4158 = (operation_194_4159);
    assign operation_194_4160 = (operation_194_4161);
    assign operation_194_4162 = ({(operation_194_4218[7:0])});
    assign operation_194_4163 = ({(operation_194_4216[7:0])});
    assign operation_194_4164 = ({(operation_194_4235[7:0])});
    assign operation_194_4165 = ({(operation_194_4189[7:0])});
    assign operation_194_4166 = ({(operation_194_4187[7:0])});
    assign operation_194_4171 = (operation_194_4172);
    assign operation_194_4173 = (operation_194_4174);
    assign operation_194_4175 = (operation_194_4176);
    assign operation_194_4177 = (operation_194_4178);
    assign operation_194_4179 = (operation_194_4180);
    assign operation_194_4181 = (operation_194_4182);
    assign operation_194_4183 = (operation_194_4184);
    assign operation_194_4185 = (operation_194_4186);
    assign operation_194_4187 = (operation_194_4188);
    assign operation_194_4189 = (operation_194_4190);
    assign operation_194_4191 = (operation_194_4192);
    assign operation_194_4199 = ({(operation_194_4234[7:0])});
    assign operation_194_4206 = ({(operation_194_4245[7:0])});
    assign operation_194_4207 = ({(operation_194_4248[7:0])});
    assign operation_194_4208 = ({(operation_194_4247[7:0])});
    assign operation_194_4209 = ({(operation_194_4250[7:0])});
    assign operation_194_4210 = ({(operation_194_4249[7:0])});
    assign operation_194_4211 = ({(operation_194_4244[7:0])});
    assign operation_194_4212 = ({(operation_194_4251[7:0])});
    assign operation_194_4213 = ({(operation_194_4246[7:0])});
    assign operation_194_4216 = (operation_194_4217);
    assign operation_194_4218 = (operation_194_4219);
    assign operation_194_4230 = ({(operation_194_4261[7:0])});
    assign operation_194_4232 = ({(operation_194_4260[7:0])});
    assign operation_194_4234 = ((control_194_27)?(lookup_sbox_31_output):(operation_194_4234_latch));
    assign operation_194_4235 = ((control_194_27)?(lookup_sbox_30_output):(operation_194_4235_latch));
    assign operation_194_4236 = ({(operation_194_4257[7:0])});
    assign operation_194_4237 = ({(operation_194_4252[7:0])});
    assign operation_194_4238 = ({(operation_194_4255[7:0])});
    assign operation_194_4239 = ({(operation_194_4258[7:0])});
    assign operation_194_4240 = ({(operation_194_4253[7:0])});
    assign operation_194_4241 = ({(operation_194_4256[7:0])});
    assign operation_194_4242 = ({(operation_194_4259[7:0])});
    assign operation_194_4243 = ({(operation_194_4254[7:0])});
    assign operation_194_4244 = ((control_194_47)?(lookup_sbox_31_output):(operation_194_4244_latch));
    assign operation_194_4245 = ((control_194_47)?(lookup_sbox_30_output):(operation_194_4245_latch));
    assign operation_194_4246 = ((control_194_47)?(lookup_sbox_29_output):(operation_194_4246_latch));
    assign operation_194_4247 = ((control_194_47)?(lookup_sbox_28_output):(operation_194_4247_latch));
    assign operation_194_4248 = ((control_194_47)?(lookup_sbox_27_output):(operation_194_4248_latch));
    assign operation_194_4249 = ((control_194_47)?(lookup_sbox_26_output):(operation_194_4249_latch));
    assign operation_194_4250 = ((control_194_47)?(lookup_sbox_25_output):(operation_194_4250_latch));
    assign operation_194_4251 = ((control_194_47)?(lookup_sbox_24_output):(operation_194_4251_latch));
    assign operation_194_4252 = ((control_194_47)?(lookup_sbox_23_output):(operation_194_4252_latch));
    assign operation_194_4253 = ((control_194_47)?(lookup_sbox_22_output):(operation_194_4253_latch));
    assign operation_194_4254 = ((control_194_47)?(lookup_sbox_21_output):(operation_194_4254_latch));
    assign operation_194_4255 = ((control_194_47)?(lookup_sbox_20_output):(operation_194_4255_latch));
    assign operation_194_4256 = ((control_194_47)?(lookup_sbox_19_output):(operation_194_4256_latch));
    assign operation_194_4257 = ((control_194_47)?(lookup_sbox_18_output):(operation_194_4257_latch));
    assign operation_194_4258 = ((control_194_47)?(lookup_sbox_17_output):(operation_194_4258_latch));
    assign operation_194_4259 = ((control_194_47)?(lookup_sbox_16_output):(operation_194_4259_latch));
    assign operation_194_4260 = ((control_194_27)?(lookup_sbox_29_output):(operation_194_4260_latch));
    assign operation_194_4261 = ((control_194_28)?(lookup_sbox_31_output):(operation_194_4261_latch));
    assign operation_194_3415 = (operation_194_3416);
    assign operation_194_3417 = ({(operation_194_3419[7:0])});
    assign operation_194_3419 = (operation_194_3420);
    assign operation_194_3421 = (operation_194_3422);
    assign operation_194_3423 = (operation_194_3424);
    assign operation_194_3425 = (operation_194_3426);
    assign operation_194_3427 = (operation_194_3428);
    assign operation_194_3429 = (operation_194_3430);
    assign operation_194_3431 = (operation_194_3432);
    assign operation_194_3433 = (operation_194_3434);
    assign operation_194_3435 = ({(operation_194_3513[7:0])});
    assign operation_194_3436 = ({(operation_194_3459[7:0])});
    assign operation_194_3437 = ({(operation_194_3457[7:0])});
    assign operation_194_3438 = ({(operation_194_3455[7:0])});
    assign operation_194_3439 = ({(operation_194_3453[7:0])});
    assign operation_194_3440 = ({(operation_194_3451[7:0])});
    assign operation_194_3441 = ({(operation_194_3449[7:0])});
    assign operation_194_3442 = ({(operation_194_3447[7:0])});
    assign operation_194_3443 = ({(operation_194_3445[7:0])});
    assign operation_194_3444 = ({(operation_194_3511[7:0])});
    assign operation_194_3445 = (operation_194_3446);
    assign operation_194_3447 = (operation_194_3448);
    assign operation_194_3449 = (operation_194_3450);
    assign operation_194_3451 = (operation_194_3452);
    assign operation_194_3453 = (operation_194_3454);
    assign operation_194_3455 = (operation_194_3456);
    assign operation_194_3457 = (operation_194_3458);
    assign operation_194_3459 = (operation_194_3460);
    assign operation_194_3461 = (operation_194_3462);
    assign operation_194_3463 = (operation_194_3464);
    assign operation_194_3465 = (operation_194_3466);
    assign operation_194_3467 = (operation_194_3468);
    assign operation_194_3469 = (operation_194_3470);
    assign operation_194_3471 = (operation_194_3472);
    assign operation_194_3473 = (operation_194_3474);
    assign operation_194_3475 = (operation_194_3476);
    assign operation_194_3477 = ({(operation_194_3543[7:0])});
    assign operation_194_3478 = ({(operation_194_3509[7:0])});
    assign operation_194_3479 = ({(operation_194_3541[7:0])});
    assign operation_194_3480 = ({(operation_194_3507[7:0])});
    assign operation_194_3481 = ({(operation_194_3505[7:0])});
    assign operation_194_3482 = ({(operation_194_3503[7:0])});
    assign operation_194_3483 = ({(operation_194_3501[7:0])});
    assign operation_194_3484 = ({(operation_194_3499[7:0])});
    assign operation_194_3485 = ({(operation_194_3497[7:0])});
    assign operation_194_3486 = ({(operation_194_3495[7:0])});
    assign operation_194_3487 = ({(operation_194_3539[7:0])});
    assign operation_194_3488 = ({(operation_194_3537[7:0])});
    assign operation_194_3489 = ({(operation_194_3535[7:0])});
    assign operation_194_3490 = ({(operation_194_3533[7:0])});
    assign operation_194_3491 = ({(operation_194_3531[7:0])});
    assign operation_194_3492 = ({(operation_194_3529[7:0])});
    assign operation_194_3493 = ({(operation_194_3527[7:0])});
    assign operation_194_3494 = ({(operation_194_3525[7:0])});
    assign operation_194_3495 = (operation_194_3496);
    assign operation_194_3497 = (operation_194_3498);
    assign operation_194_3499 = (operation_194_3500);
    assign operation_194_3501 = (operation_194_3502);
    assign operation_194_3503 = (operation_194_3504);
    assign operation_194_3505 = (operation_194_3506);
    assign operation_194_3507 = (operation_194_3508);
    assign operation_194_3509 = (operation_194_3510);
    assign operation_194_3511 = (operation_194_3512);
    assign operation_194_3513 = (operation_194_3514);
    assign operation_194_3515 = ({(operation_194_3573[7:0])});
    assign operation_194_3516 = ({(operation_194_3571[7:0])});
    assign operation_194_3517 = ({(operation_194_3569[7:0])});
    assign operation_194_3518 = ({(operation_194_3567[7:0])});
    assign operation_194_3519 = ({(operation_194_3565[7:0])});
    assign operation_194_3520 = ({(operation_194_3563[7:0])});
    assign operation_194_3521 = ({(operation_194_3561[7:0])});
    assign operation_194_3522 = ({(operation_194_3559[7:0])});
    assign operation_194_3523 = ({(operation_194_3557[7:0])});
    assign operation_194_3524 = ({(operation_194_3555[7:0])});
    assign operation_194_3525 = (operation_194_3526);
    assign operation_194_3527 = (operation_194_3528);
    assign operation_194_3529 = (operation_194_3530);
    assign operation_194_3531 = (operation_194_3532);
    assign operation_194_3533 = (operation_194_3534);
    assign operation_194_3535 = (operation_194_3536);
    assign operation_194_3537 = (operation_194_3538);
    assign operation_194_3539 = (operation_194_3540);
    assign operation_194_3541 = (operation_194_3542);
    assign operation_194_3543 = (operation_194_3544);
    assign operation_194_3545 = ({(operation_194_3611[7:0])});
    assign operation_194_3546 = ({(operation_194_3609[7:0])});
    assign operation_194_3547 = ({(operation_194_3606[7:0])});
    assign operation_194_3548 = ({(operation_194_3603[7:0])});
    assign operation_194_3549 = ({(operation_194_3600[7:0])});
    assign operation_194_3550 = ({(operation_194_3597[7:0])});
    assign operation_194_3551 = ({(operation_194_3594[7:0])});
    assign operation_194_3552 = ({(operation_194_3591[7:0])});
    assign operation_194_3553 = ({(operation_194_3588[7:0])});
    assign operation_194_3554 = ({(operation_194_3585[7:0])});
    assign operation_194_3555 = (operation_194_3556);
    assign operation_194_3557 = (operation_194_3558);
    assign operation_194_3559 = (operation_194_3560);
    assign operation_194_3561 = (operation_194_3562);
    assign operation_194_3563 = (operation_194_3564);
    assign operation_194_3565 = (operation_194_3566);
    assign operation_194_3567 = (operation_194_3568);
    assign operation_194_3569 = (operation_194_3570);
    assign operation_194_3571 = (operation_194_3572);
    assign operation_194_3573 = (operation_194_3574);
    assign operation_194_3575 = ({(operation_194_3673[7:0])});
    assign operation_194_3576 = ({(operation_194_3671[7:0])});
    assign operation_194_3577 = ({(operation_194_3668[7:0])});
    assign operation_194_3578 = ({(operation_194_3665[7:0])});
    assign operation_194_3579 = ({(operation_194_3662[7:0])});
    assign operation_194_3580 = ({(operation_194_3659[7:0])});
    assign operation_194_3581 = ({(operation_194_3656[7:0])});
    assign operation_194_3582 = ({(operation_194_3653[7:0])});
    assign operation_194_3583 = ({(operation_194_3650[7:0])});
    assign operation_194_3584 = ({(operation_194_3647[7:0])});
    assign operation_194_3585 = (operation_194_3586);
    assign operation_194_3588 = (operation_194_3589);
    assign operation_194_3591 = (operation_194_3592);
    assign operation_194_3594 = (operation_194_3595);
    assign operation_194_3597 = (operation_194_3598);
    assign operation_194_3600 = (operation_194_3601);
    assign operation_194_3603 = (operation_194_3604);
    assign operation_194_3606 = (operation_194_3607);
    assign operation_194_3609 = (operation_194_3610);
    assign operation_194_3611 = (operation_194_3612);
    assign operation_194_3613 = ({(operation_194_3731[7:0])});
    assign operation_194_3614 = ({(operation_194_3729[7:0])});
    assign operation_194_3618 = ({(operation_194_3721[7:0])});
    assign operation_194_3622 = ({(operation_194_3720[7:0])});
    assign operation_194_3626 = ({(operation_194_3718[7:0])});
    assign operation_194_3630 = ({(operation_194_3717[7:0])});
    assign operation_194_3634 = ({(operation_194_3715[7:0])});
    assign operation_194_3638 = ({(operation_194_3714[7:0])});
    assign operation_194_3642 = ({(operation_194_3712[7:0])});
    assign operation_194_3646 = ({(operation_194_3711[7:0])});
    assign operation_194_3647 = (operation_194_3648);
    assign operation_194_3650 = (operation_194_3651);
    assign operation_194_3653 = (operation_194_3654);
    assign operation_194_3656 = (operation_194_3657);
    assign operation_194_3659 = (operation_194_3660);
    assign operation_194_3662 = (operation_194_3663);
    assign operation_194_3665 = (operation_194_3666);
    assign operation_194_3668 = (operation_194_3669);
    assign operation_194_3671 = (operation_194_3672);
    assign operation_194_3673 = (operation_194_3674);
    assign operation_194_3675 = ({(operation_194_3762[7:0])});
    assign operation_194_3676 = ({(operation_194_3727[7:0])});
    assign operation_194_3677 = ({(operation_194_3725[7:0])});
    assign operation_194_3678 = ({(operation_194_3723[7:0])});
    assign operation_194_3682 = ({(operation_194_3756[7:0])});
    assign operation_194_3686 = ({(operation_194_3754[7:0])});
    assign operation_194_3690 = ({(operation_194_3752[7:0])});
    assign operation_194_3694 = ({(operation_194_3750[7:0])});
    assign operation_194_3698 = ({(operation_194_3748[7:0])});
    assign operation_194_3702 = ({(operation_194_3746[7:0])});
    assign operation_194_3706 = ({(operation_194_3744[7:0])});
    assign operation_194_3710 = ({(operation_194_3742[7:0])});
    assign operation_194_3711 = (operation_194_3741);
    assign operation_194_3712 = (operation_194_3713);
    assign operation_194_3714 = (operation_194_3776);
    assign operation_194_3715 = (operation_194_3716);
    assign operation_194_3717 = (operation_194_3739);
    assign operation_194_3718 = (operation_194_3719);
    assign operation_194_3720 = (operation_194_3774);
    assign operation_194_3721 = (operation_194_3722);
    assign operation_194_3723 = (operation_194_3724);
    assign operation_194_3725 = (operation_194_3726);
    assign operation_194_3727 = (operation_194_3728);
    assign operation_194_3729 = (operation_194_3730);
    assign operation_194_3731 = (operation_194_3732);
    assign operation_194_3733 = ({(operation_194_3789[7:0])});
    assign operation_194_3734 = ({(operation_194_3787[7:0])});
    assign operation_194_3735 = ({(operation_194_3806[7:0])});
    assign operation_194_3736 = ({(operation_194_3760[7:0])});
    assign operation_194_3737 = ({(operation_194_3758[7:0])});
    assign operation_194_3742 = (operation_194_3743);
    assign operation_194_3744 = (operation_194_3745);
    assign operation_194_3746 = (operation_194_3747);
    assign operation_194_3748 = (operation_194_3749);
    assign operation_194_3750 = (operation_194_3751);
    assign operation_194_3752 = (operation_194_3753);
    assign operation_194_3754 = (operation_194_3755);
    assign operation_194_3756 = (operation_194_3757);
    assign operation_194_3758 = (operation_194_3759);
    assign operation_194_3760 = (operation_194_3761);
    assign operation_194_3762 = (operation_194_3763);
    assign operation_194_3770 = ({(operation_194_3805[7:0])});
    assign operation_194_3777 = ({(operation_194_3816[7:0])});
    assign operation_194_3778 = ({(operation_194_3819[7:0])});
    assign operation_194_3779 = ({(operation_194_3818[7:0])});
    assign operation_194_3780 = ({(operation_194_3821[7:0])});
    assign operation_194_3781 = ({(operation_194_3820[7:0])});
    assign operation_194_3782 = ({(operation_194_3815[7:0])});
    assign operation_194_3783 = ({(operation_194_3822[7:0])});
    assign operation_194_3784 = ({(operation_194_3817[7:0])});
    assign operation_194_3787 = (operation_194_3788);
    assign operation_194_3789 = (operation_194_3790);
    assign operation_194_3801 = ({(operation_194_3832[7:0])});
    assign operation_194_3803 = ({(operation_194_3831[7:0])});
    assign operation_194_3805 = ((control_194_22)?(lookup_sbox_31_output):(operation_194_3805_latch));
    assign operation_194_3806 = ((control_194_22)?(lookup_sbox_30_output):(operation_194_3806_latch));
    assign operation_194_3807 = ({(operation_194_3828[7:0])});
    assign operation_194_3808 = ({(operation_194_3823[7:0])});
    assign operation_194_3809 = ({(operation_194_3826[7:0])});
    assign operation_194_3810 = ({(operation_194_3829[7:0])});
    assign operation_194_3811 = ({(operation_194_3824[7:0])});
    assign operation_194_3812 = ({(operation_194_3827[7:0])});
    assign operation_194_3813 = ({(operation_194_3830[7:0])});
    assign operation_194_3814 = ({(operation_194_3825[7:0])});
    assign operation_194_3815 = ((control_194_38)?(lookup_sbox_28_output):(operation_194_3815_latch));
    assign operation_194_3816 = ((control_194_38)?(lookup_sbox_27_output):(operation_194_3816_latch));
    assign operation_194_3817 = ((control_194_38)?(lookup_sbox_26_output):(operation_194_3817_latch));
    assign operation_194_3818 = ((control_194_38)?(lookup_sbox_25_output):(operation_194_3818_latch));
    assign operation_194_3819 = ((control_194_38)?(lookup_sbox_24_output):(operation_194_3819_latch));
    assign operation_194_3820 = ((control_194_38)?(lookup_sbox_23_output):(operation_194_3820_latch));
    assign operation_194_3821 = ((control_194_38)?(lookup_sbox_22_output):(operation_194_3821_latch));
    assign operation_194_3822 = ((control_194_38)?(lookup_sbox_21_output):(operation_194_3822_latch));
    assign operation_194_3823 = ((control_194_38)?(lookup_sbox_20_output):(operation_194_3823_latch));
    assign operation_194_3824 = ((control_194_38)?(lookup_sbox_19_output):(operation_194_3824_latch));
    assign operation_194_3825 = ((control_194_38)?(lookup_sbox_18_output):(operation_194_3825_latch));
    assign operation_194_3826 = ((control_194_38)?(lookup_sbox_17_output):(operation_194_3826_latch));
    assign operation_194_3827 = ((control_194_38)?(lookup_sbox_16_output):(operation_194_3827_latch));
    assign operation_194_3828 = ((control_194_38)?(lookup_sbox_15_output):(operation_194_3828_latch));
    assign operation_194_3829 = ((control_194_38)?(lookup_sbox_14_output):(operation_194_3829_latch));
    assign operation_194_3830 = ((control_194_38)?(lookup_sbox_13_output):(operation_194_3830_latch));
    assign operation_194_3831 = ((control_194_22)?(lookup_sbox_29_output):(operation_194_3831_latch));
    assign operation_194_3832 = ((control_194_22)?(lookup_sbox_28_output):(operation_194_3832_latch));
    assign operation_194_2986 = (operation_194_2987);
    assign operation_194_2988 = ({(operation_194_2990[7:0])});
    assign operation_194_2990 = (operation_194_2991);
    assign operation_194_2992 = (operation_194_2993);
    assign operation_194_2994 = (operation_194_2995);
    assign operation_194_2996 = (operation_194_2997);
    assign operation_194_2998 = (operation_194_2999);
    assign operation_194_3000 = (operation_194_3001);
    assign operation_194_3002 = (operation_194_3003);
    assign operation_194_3004 = (operation_194_3005);
    assign operation_194_3006 = ({(operation_194_3084[7:0])});
    assign operation_194_3007 = ({(operation_194_3030[7:0])});
    assign operation_194_3008 = ({(operation_194_3028[7:0])});
    assign operation_194_3009 = ({(operation_194_3026[7:0])});
    assign operation_194_3010 = ({(operation_194_3024[7:0])});
    assign operation_194_3011 = ({(operation_194_3022[7:0])});
    assign operation_194_3012 = ({(operation_194_3020[7:0])});
    assign operation_194_3013 = ({(operation_194_3018[7:0])});
    assign operation_194_3014 = ({(operation_194_3016[7:0])});
    assign operation_194_3015 = ({(operation_194_3082[7:0])});
    assign operation_194_3016 = (operation_194_3017);
    assign operation_194_3018 = (operation_194_3019);
    assign operation_194_3020 = (operation_194_3021);
    assign operation_194_3022 = (operation_194_3023);
    assign operation_194_3024 = (operation_194_3025);
    assign operation_194_3026 = (operation_194_3027);
    assign operation_194_3028 = (operation_194_3029);
    assign operation_194_3030 = (operation_194_3031);
    assign operation_194_3032 = (operation_194_3033);
    assign operation_194_3034 = (operation_194_3035);
    assign operation_194_3036 = (operation_194_3037);
    assign operation_194_3038 = (operation_194_3039);
    assign operation_194_3040 = (operation_194_3041);
    assign operation_194_3042 = (operation_194_3043);
    assign operation_194_3044 = (operation_194_3045);
    assign operation_194_3046 = (operation_194_3047);
    assign operation_194_3048 = ({(operation_194_3114[7:0])});
    assign operation_194_3049 = ({(operation_194_3080[7:0])});
    assign operation_194_3050 = ({(operation_194_3112[7:0])});
    assign operation_194_3051 = ({(operation_194_3078[7:0])});
    assign operation_194_3052 = ({(operation_194_3076[7:0])});
    assign operation_194_3053 = ({(operation_194_3074[7:0])});
    assign operation_194_3054 = ({(operation_194_3072[7:0])});
    assign operation_194_3055 = ({(operation_194_3070[7:0])});
    assign operation_194_3056 = ({(operation_194_3068[7:0])});
    assign operation_194_3057 = ({(operation_194_3066[7:0])});
    assign operation_194_3058 = ({(operation_194_3110[7:0])});
    assign operation_194_3059 = ({(operation_194_3108[7:0])});
    assign operation_194_3060 = ({(operation_194_3106[7:0])});
    assign operation_194_3061 = ({(operation_194_3104[7:0])});
    assign operation_194_3062 = ({(operation_194_3102[7:0])});
    assign operation_194_3063 = ({(operation_194_3100[7:0])});
    assign operation_194_3064 = ({(operation_194_3098[7:0])});
    assign operation_194_3065 = ({(operation_194_3096[7:0])});
    assign operation_194_3066 = (operation_194_3067);
    assign operation_194_3068 = (operation_194_3069);
    assign operation_194_3070 = (operation_194_3071);
    assign operation_194_3072 = (operation_194_3073);
    assign operation_194_3074 = (operation_194_3075);
    assign operation_194_3076 = (operation_194_3077);
    assign operation_194_3078 = (operation_194_3079);
    assign operation_194_3080 = (operation_194_3081);
    assign operation_194_3082 = (operation_194_3083);
    assign operation_194_3084 = (operation_194_3085);
    assign operation_194_3086 = ({(operation_194_3144[7:0])});
    assign operation_194_3087 = ({(operation_194_3142[7:0])});
    assign operation_194_3088 = ({(operation_194_3140[7:0])});
    assign operation_194_3089 = ({(operation_194_3138[7:0])});
    assign operation_194_3090 = ({(operation_194_3136[7:0])});
    assign operation_194_3091 = ({(operation_194_3134[7:0])});
    assign operation_194_3092 = ({(operation_194_3132[7:0])});
    assign operation_194_3093 = ({(operation_194_3130[7:0])});
    assign operation_194_3094 = ({(operation_194_3128[7:0])});
    assign operation_194_3095 = ({(operation_194_3126[7:0])});
    assign operation_194_3096 = (operation_194_3097);
    assign operation_194_3098 = (operation_194_3099);
    assign operation_194_3100 = (operation_194_3101);
    assign operation_194_3102 = (operation_194_3103);
    assign operation_194_3104 = (operation_194_3105);
    assign operation_194_3106 = (operation_194_3107);
    assign operation_194_3108 = (operation_194_3109);
    assign operation_194_3110 = (operation_194_3111);
    assign operation_194_3112 = (operation_194_3113);
    assign operation_194_3114 = (operation_194_3115);
    assign operation_194_3116 = ({(operation_194_3182[7:0])});
    assign operation_194_3117 = ({(operation_194_3180[7:0])});
    assign operation_194_3118 = ({(operation_194_3177[7:0])});
    assign operation_194_3119 = ({(operation_194_3174[7:0])});
    assign operation_194_3120 = ({(operation_194_3171[7:0])});
    assign operation_194_3121 = ({(operation_194_3168[7:0])});
    assign operation_194_3122 = ({(operation_194_3165[7:0])});
    assign operation_194_3123 = ({(operation_194_3162[7:0])});
    assign operation_194_3124 = ({(operation_194_3159[7:0])});
    assign operation_194_3125 = ({(operation_194_3156[7:0])});
    assign operation_194_3126 = (operation_194_3127);
    assign operation_194_3128 = (operation_194_3129);
    assign operation_194_3130 = (operation_194_3131);
    assign operation_194_3132 = (operation_194_3133);
    assign operation_194_3134 = (operation_194_3135);
    assign operation_194_3136 = (operation_194_3137);
    assign operation_194_3138 = (operation_194_3139);
    assign operation_194_3140 = (operation_194_3141);
    assign operation_194_3142 = (operation_194_3143);
    assign operation_194_3144 = (operation_194_3145);
    assign operation_194_3146 = ({(operation_194_3244[7:0])});
    assign operation_194_3147 = ({(operation_194_3242[7:0])});
    assign operation_194_3148 = ({(operation_194_3239[7:0])});
    assign operation_194_3149 = ({(operation_194_3236[7:0])});
    assign operation_194_3150 = ({(operation_194_3233[7:0])});
    assign operation_194_3151 = ({(operation_194_3230[7:0])});
    assign operation_194_3152 = ({(operation_194_3227[7:0])});
    assign operation_194_3153 = ({(operation_194_3224[7:0])});
    assign operation_194_3154 = ({(operation_194_3221[7:0])});
    assign operation_194_3155 = ({(operation_194_3218[7:0])});
    assign operation_194_3156 = (operation_194_3157);
    assign operation_194_3159 = (operation_194_3160);
    assign operation_194_3162 = (operation_194_3163);
    assign operation_194_3165 = (operation_194_3166);
    assign operation_194_3168 = (operation_194_3169);
    assign operation_194_3171 = (operation_194_3172);
    assign operation_194_3174 = (operation_194_3175);
    assign operation_194_3177 = (operation_194_3178);
    assign operation_194_3180 = (operation_194_3181);
    assign operation_194_3182 = (operation_194_3183);
    assign operation_194_3184 = ({(operation_194_3302[7:0])});
    assign operation_194_3185 = ({(operation_194_3300[7:0])});
    assign operation_194_3189 = ({(operation_194_3292[7:0])});
    assign operation_194_3193 = ({(operation_194_3291[7:0])});
    assign operation_194_3197 = ({(operation_194_3289[7:0])});
    assign operation_194_3201 = ({(operation_194_3288[7:0])});
    assign operation_194_3205 = ({(operation_194_3286[7:0])});
    assign operation_194_3209 = ({(operation_194_3285[7:0])});
    assign operation_194_3213 = ({(operation_194_3283[7:0])});
    assign operation_194_3217 = ({(operation_194_3282[7:0])});
    assign operation_194_3218 = (operation_194_3219);
    assign operation_194_3221 = (operation_194_3222);
    assign operation_194_3224 = (operation_194_3225);
    assign operation_194_3227 = (operation_194_3228);
    assign operation_194_3230 = (operation_194_3231);
    assign operation_194_3233 = (operation_194_3234);
    assign operation_194_3236 = (operation_194_3237);
    assign operation_194_3239 = (operation_194_3240);
    assign operation_194_3242 = (operation_194_3243);
    assign operation_194_3244 = (operation_194_3245);
    assign operation_194_3246 = ({(operation_194_3333[7:0])});
    assign operation_194_3247 = ({(operation_194_3298[7:0])});
    assign operation_194_3248 = ({(operation_194_3296[7:0])});
    assign operation_194_3249 = ({(operation_194_3294[7:0])});
    assign operation_194_3253 = ({(operation_194_3327[7:0])});
    assign operation_194_3257 = ({(operation_194_3325[7:0])});
    assign operation_194_3261 = ({(operation_194_3323[7:0])});
    assign operation_194_3265 = ({(operation_194_3321[7:0])});
    assign operation_194_3269 = ({(operation_194_3319[7:0])});
    assign operation_194_3273 = ({(operation_194_3317[7:0])});
    assign operation_194_3277 = ({(operation_194_3315[7:0])});
    assign operation_194_3281 = ({(operation_194_3313[7:0])});
    assign operation_194_3282 = (operation_194_3312);
    assign operation_194_3283 = (operation_194_3284);
    assign operation_194_3285 = (operation_194_3347);
    assign operation_194_3286 = (operation_194_3287);
    assign operation_194_3288 = (operation_194_3310);
    assign operation_194_3289 = (operation_194_3290);
    assign operation_194_3291 = (operation_194_3345);
    assign operation_194_3292 = (operation_194_3293);
    assign operation_194_3294 = (operation_194_3295);
    assign operation_194_3296 = (operation_194_3297);
    assign operation_194_3298 = (operation_194_3299);
    assign operation_194_3300 = (operation_194_3301);
    assign operation_194_3302 = (operation_194_3303);
    assign operation_194_3304 = ({(operation_194_3360[7:0])});
    assign operation_194_3305 = ({(operation_194_3358[7:0])});
    assign operation_194_3306 = ({(operation_194_3377[7:0])});
    assign operation_194_3307 = ({(operation_194_3331[7:0])});
    assign operation_194_3308 = ({(operation_194_3329[7:0])});
    assign operation_194_3313 = (operation_194_3314);
    assign operation_194_3315 = (operation_194_3316);
    assign operation_194_3317 = (operation_194_3318);
    assign operation_194_3319 = (operation_194_3320);
    assign operation_194_3321 = (operation_194_3322);
    assign operation_194_3323 = (operation_194_3324);
    assign operation_194_3325 = (operation_194_3326);
    assign operation_194_3327 = (operation_194_3328);
    assign operation_194_3329 = (operation_194_3330);
    assign operation_194_3331 = (operation_194_3332);
    assign operation_194_3333 = (operation_194_3334);
    assign operation_194_3341 = ({(operation_194_3376[7:0])});
    assign operation_194_3348 = ({(operation_194_3387[7:0])});
    assign operation_194_3349 = ({(operation_194_3390[7:0])});
    assign operation_194_3350 = ({(operation_194_3389[7:0])});
    assign operation_194_3351 = ({(operation_194_3392[7:0])});
    assign operation_194_3352 = ({(operation_194_3391[7:0])});
    assign operation_194_3353 = ({(operation_194_3386[7:0])});
    assign operation_194_3354 = ({(operation_194_3393[7:0])});
    assign operation_194_3355 = ({(operation_194_3388[7:0])});
    assign operation_194_3358 = (operation_194_3359);
    assign operation_194_3360 = (operation_194_3361);
    assign operation_194_3372 = ({(operation_194_3403[7:0])});
    assign operation_194_3374 = ({(operation_194_3402[7:0])});
    assign operation_194_3376 = ((control_194_17)?(lookup_sbox_31_output):(operation_194_3376_latch));
    assign operation_194_3377 = ((control_194_16)?(lookup_sbox_31_output):(operation_194_3377_latch));
    assign operation_194_3378 = ({(operation_194_3399[7:0])});
    assign operation_194_3379 = ({(operation_194_3394[7:0])});
    assign operation_194_3380 = ({(operation_194_3397[7:0])});
    assign operation_194_3381 = ({(operation_194_3400[7:0])});
    assign operation_194_3382 = ({(operation_194_3395[7:0])});
    assign operation_194_3383 = ({(operation_194_3398[7:0])});
    assign operation_194_3384 = ({(operation_194_3401[7:0])});
    assign operation_194_3385 = ({(operation_194_3396[7:0])});
    assign operation_194_3386 = ((control_194_29)?(lookup_sbox_31_output):(operation_194_3386_latch));
    assign operation_194_3387 = ((control_194_29)?(lookup_sbox_30_output):(operation_194_3387_latch));
    assign operation_194_3388 = ((control_194_29)?(lookup_sbox_29_output):(operation_194_3388_latch));
    assign operation_194_3389 = ((control_194_29)?(lookup_sbox_28_output):(operation_194_3389_latch));
    assign operation_194_3390 = ((control_194_29)?(lookup_sbox_27_output):(operation_194_3390_latch));
    assign operation_194_3391 = ((control_194_29)?(lookup_sbox_26_output):(operation_194_3391_latch));
    assign operation_194_3392 = ((control_194_29)?(lookup_sbox_25_output):(operation_194_3392_latch));
    assign operation_194_3393 = ((control_194_29)?(lookup_sbox_24_output):(operation_194_3393_latch));
    assign operation_194_3394 = ((control_194_29)?(lookup_sbox_23_output):(operation_194_3394_latch));
    assign operation_194_3395 = ((control_194_29)?(lookup_sbox_22_output):(operation_194_3395_latch));
    assign operation_194_3396 = ((control_194_29)?(lookup_sbox_21_output):(operation_194_3396_latch));
    assign operation_194_3397 = ((control_194_29)?(lookup_sbox_20_output):(operation_194_3397_latch));
    assign operation_194_3398 = ((control_194_29)?(lookup_sbox_19_output):(operation_194_3398_latch));
    assign operation_194_3399 = ((control_194_29)?(lookup_sbox_18_output):(operation_194_3399_latch));
    assign operation_194_3400 = ((control_194_29)?(lookup_sbox_17_output):(operation_194_3400_latch));
    assign operation_194_3401 = ((control_194_29)?(lookup_sbox_16_output):(operation_194_3401_latch));
    assign operation_194_3402 = ((control_194_17)?(lookup_sbox_30_output):(operation_194_3402_latch));
    assign operation_194_3403 = ((control_194_17)?(lookup_sbox_29_output):(operation_194_3403_latch));
    assign operation_194_2557 = (operation_194_2558);
    assign operation_194_2559 = ({(operation_194_2561[7:0])});
    assign operation_194_2561 = (operation_194_2562);
    assign operation_194_2563 = (operation_194_2564);
    assign operation_194_2565 = (operation_194_2566);
    assign operation_194_2567 = (operation_194_2568);
    assign operation_194_2569 = (operation_194_2570);
    assign operation_194_2571 = (operation_194_2572);
    assign operation_194_2573 = (operation_194_2574);
    assign operation_194_2575 = (operation_194_2576);
    assign operation_194_2577 = ({(operation_194_2655[7:0])});
    assign operation_194_2578 = ({(operation_194_2601[7:0])});
    assign operation_194_2579 = ({(operation_194_2599[7:0])});
    assign operation_194_2580 = ({(operation_194_2597[7:0])});
    assign operation_194_2581 = ({(operation_194_2595[7:0])});
    assign operation_194_2582 = ({(operation_194_2593[7:0])});
    assign operation_194_2583 = ({(operation_194_2591[7:0])});
    assign operation_194_2584 = ({(operation_194_2589[7:0])});
    assign operation_194_2585 = ({(operation_194_2587[7:0])});
    assign operation_194_2586 = ({(operation_194_2653[7:0])});
    assign operation_194_2587 = (operation_194_2588);
    assign operation_194_2589 = (operation_194_2590);
    assign operation_194_2591 = (operation_194_2592);
    assign operation_194_2593 = (operation_194_2594);
    assign operation_194_2595 = (operation_194_2596);
    assign operation_194_2597 = (operation_194_2598);
    assign operation_194_2599 = (operation_194_2600);
    assign operation_194_2601 = (operation_194_2602);
    assign operation_194_2603 = (operation_194_2604);
    assign operation_194_2605 = (operation_194_2606);
    assign operation_194_2607 = (operation_194_2608);
    assign operation_194_2609 = (operation_194_2610);
    assign operation_194_2611 = (operation_194_2612);
    assign operation_194_2613 = (operation_194_2614);
    assign operation_194_2615 = (operation_194_2616);
    assign operation_194_2617 = (operation_194_2618);
    assign operation_194_2619 = ({(operation_194_2685[7:0])});
    assign operation_194_2620 = ({(operation_194_2651[7:0])});
    assign operation_194_2621 = ({(operation_194_2683[7:0])});
    assign operation_194_2622 = ({(operation_194_2649[7:0])});
    assign operation_194_2623 = ({(operation_194_2647[7:0])});
    assign operation_194_2624 = ({(operation_194_2645[7:0])});
    assign operation_194_2625 = ({(operation_194_2643[7:0])});
    assign operation_194_2626 = ({(operation_194_2641[7:0])});
    assign operation_194_2627 = ({(operation_194_2639[7:0])});
    assign operation_194_2628 = ({(operation_194_2637[7:0])});
    assign operation_194_2629 = ({(operation_194_2681[7:0])});
    assign operation_194_2630 = ({(operation_194_2679[7:0])});
    assign operation_194_2631 = ({(operation_194_2677[7:0])});
    assign operation_194_2632 = ({(operation_194_2675[7:0])});
    assign operation_194_2633 = ({(operation_194_2673[7:0])});
    assign operation_194_2634 = ({(operation_194_2671[7:0])});
    assign operation_194_2635 = ({(operation_194_2669[7:0])});
    assign operation_194_2636 = ({(operation_194_2667[7:0])});
    assign operation_194_2637 = (operation_194_2638);
    assign operation_194_2639 = (operation_194_2640);
    assign operation_194_2641 = (operation_194_2642);
    assign operation_194_2643 = (operation_194_2644);
    assign operation_194_2645 = (operation_194_2646);
    assign operation_194_2647 = (operation_194_2648);
    assign operation_194_2649 = (operation_194_2650);
    assign operation_194_2651 = (operation_194_2652);
    assign operation_194_2653 = (operation_194_2654);
    assign operation_194_2655 = (operation_194_2656);
    assign operation_194_2657 = ({(operation_194_2715[7:0])});
    assign operation_194_2658 = ({(operation_194_2713[7:0])});
    assign operation_194_2659 = ({(operation_194_2711[7:0])});
    assign operation_194_2660 = ({(operation_194_2709[7:0])});
    assign operation_194_2661 = ({(operation_194_2707[7:0])});
    assign operation_194_2662 = ({(operation_194_2705[7:0])});
    assign operation_194_2663 = ({(operation_194_2703[7:0])});
    assign operation_194_2664 = ({(operation_194_2701[7:0])});
    assign operation_194_2665 = ({(operation_194_2699[7:0])});
    assign operation_194_2666 = ({(operation_194_2697[7:0])});
    assign operation_194_2667 = (operation_194_2668);
    assign operation_194_2669 = (operation_194_2670);
    assign operation_194_2671 = (operation_194_2672);
    assign operation_194_2673 = (operation_194_2674);
    assign operation_194_2675 = (operation_194_2676);
    assign operation_194_2677 = (operation_194_2678);
    assign operation_194_2679 = (operation_194_2680);
    assign operation_194_2681 = (operation_194_2682);
    assign operation_194_2683 = (operation_194_2684);
    assign operation_194_2685 = (operation_194_2686);
    assign operation_194_2687 = ({(operation_194_2753[7:0])});
    assign operation_194_2688 = ({(operation_194_2751[7:0])});
    assign operation_194_2689 = ({(operation_194_2748[7:0])});
    assign operation_194_2690 = ({(operation_194_2745[7:0])});
    assign operation_194_2691 = ({(operation_194_2742[7:0])});
    assign operation_194_2692 = ({(operation_194_2739[7:0])});
    assign operation_194_2693 = ({(operation_194_2736[7:0])});
    assign operation_194_2694 = ({(operation_194_2733[7:0])});
    assign operation_194_2695 = ({(operation_194_2730[7:0])});
    assign operation_194_2696 = ({(operation_194_2727[7:0])});
    assign operation_194_2697 = (operation_194_2698);
    assign operation_194_2699 = (operation_194_2700);
    assign operation_194_2701 = (operation_194_2702);
    assign operation_194_2703 = (operation_194_2704);
    assign operation_194_2705 = (operation_194_2706);
    assign operation_194_2707 = (operation_194_2708);
    assign operation_194_2709 = (operation_194_2710);
    assign operation_194_2711 = (operation_194_2712);
    assign operation_194_2713 = (operation_194_2714);
    assign operation_194_2715 = (operation_194_2716);
    assign operation_194_2717 = ({(operation_194_2815[7:0])});
    assign operation_194_2718 = ({(operation_194_2813[7:0])});
    assign operation_194_2719 = ({(operation_194_2810[7:0])});
    assign operation_194_2720 = ({(operation_194_2807[7:0])});
    assign operation_194_2721 = ({(operation_194_2804[7:0])});
    assign operation_194_2722 = ({(operation_194_2801[7:0])});
    assign operation_194_2723 = ({(operation_194_2798[7:0])});
    assign operation_194_2724 = ({(operation_194_2795[7:0])});
    assign operation_194_2725 = ({(operation_194_2792[7:0])});
    assign operation_194_2726 = ({(operation_194_2789[7:0])});
    assign operation_194_2727 = (operation_194_2728);
    assign operation_194_2730 = (operation_194_2731);
    assign operation_194_2733 = (operation_194_2734);
    assign operation_194_2736 = (operation_194_2737);
    assign operation_194_2739 = (operation_194_2740);
    assign operation_194_2742 = (operation_194_2743);
    assign operation_194_2745 = (operation_194_2746);
    assign operation_194_2748 = (operation_194_2749);
    assign operation_194_2751 = (operation_194_2752);
    assign operation_194_2753 = (operation_194_2754);
    assign operation_194_2755 = ({(operation_194_2873[7:0])});
    assign operation_194_2756 = ({(operation_194_2871[7:0])});
    assign operation_194_2760 = ({(operation_194_2863[7:0])});
    assign operation_194_2764 = ({(operation_194_2862[7:0])});
    assign operation_194_2768 = ({(operation_194_2860[7:0])});
    assign operation_194_2772 = ({(operation_194_2859[7:0])});
    assign operation_194_2776 = ({(operation_194_2857[7:0])});
    assign operation_194_2780 = ({(operation_194_2856[7:0])});
    assign operation_194_2784 = ({(operation_194_2854[7:0])});
    assign operation_194_2788 = ({(operation_194_2853[7:0])});
    assign operation_194_2789 = (operation_194_2790);
    assign operation_194_2792 = (operation_194_2793);
    assign operation_194_2795 = (operation_194_2796);
    assign operation_194_2798 = (operation_194_2799);
    assign operation_194_2801 = (operation_194_2802);
    assign operation_194_2804 = (operation_194_2805);
    assign operation_194_2807 = (operation_194_2808);
    assign operation_194_2810 = (operation_194_2811);
    assign operation_194_2813 = (operation_194_2814);
    assign operation_194_2815 = (operation_194_2816);
    assign operation_194_2817 = ({(operation_194_2904[7:0])});
    assign operation_194_2818 = ({(operation_194_2869[7:0])});
    assign operation_194_2819 = ({(operation_194_2867[7:0])});
    assign operation_194_2820 = ({(operation_194_2865[7:0])});
    assign operation_194_2824 = ({(operation_194_2898[7:0])});
    assign operation_194_2828 = ({(operation_194_2896[7:0])});
    assign operation_194_2832 = ({(operation_194_2894[7:0])});
    assign operation_194_2836 = ({(operation_194_2892[7:0])});
    assign operation_194_2840 = ({(operation_194_2890[7:0])});
    assign operation_194_2844 = ({(operation_194_2888[7:0])});
    assign operation_194_2848 = ({(operation_194_2886[7:0])});
    assign operation_194_2852 = ({(operation_194_2884[7:0])});
    assign operation_194_2853 = (operation_194_2883);
    assign operation_194_2854 = (operation_194_2855);
    assign operation_194_2856 = (operation_194_2918);
    assign operation_194_2857 = (operation_194_2858);
    assign operation_194_2859 = (operation_194_2881);
    assign operation_194_2860 = (operation_194_2861);
    assign operation_194_2862 = (operation_194_2916);
    assign operation_194_2863 = (operation_194_2864);
    assign operation_194_2865 = (operation_194_2866);
    assign operation_194_2867 = (operation_194_2868);
    assign operation_194_2869 = (operation_194_2870);
    assign operation_194_2871 = (operation_194_2872);
    assign operation_194_2873 = (operation_194_2874);
    assign operation_194_2875 = ({(operation_194_2931[7:0])});
    assign operation_194_2876 = ({(operation_194_2929[7:0])});
    assign operation_194_2877 = ({(operation_194_2948[7:0])});
    assign operation_194_2878 = ({(operation_194_2902[7:0])});
    assign operation_194_2879 = ({(operation_194_2900[7:0])});
    assign operation_194_2884 = (operation_194_2885);
    assign operation_194_2886 = (operation_194_2887);
    assign operation_194_2888 = (operation_194_2889);
    assign operation_194_2890 = (operation_194_2891);
    assign operation_194_2892 = (operation_194_2893);
    assign operation_194_2894 = (operation_194_2895);
    assign operation_194_2896 = (operation_194_2897);
    assign operation_194_2898 = (operation_194_2899);
    assign operation_194_2900 = (operation_194_2901);
    assign operation_194_2902 = (operation_194_2903);
    assign operation_194_2904 = (operation_194_2905);
    assign operation_194_2912 = ({(operation_194_2947[7:0])});
    assign operation_194_2919 = ({(operation_194_2958[7:0])});
    assign operation_194_2920 = ({(operation_194_2961[7:0])});
    assign operation_194_2921 = ({(operation_194_2960[7:0])});
    assign operation_194_2922 = ({(operation_194_2963[7:0])});
    assign operation_194_2923 = ({(operation_194_2962[7:0])});
    assign operation_194_2924 = ({(operation_194_2957[7:0])});
    assign operation_194_2925 = ({(operation_194_2964[7:0])});
    assign operation_194_2926 = ({(operation_194_2959[7:0])});
    assign operation_194_2929 = (operation_194_2930);
    assign operation_194_2931 = (operation_194_2932);
    assign operation_194_2943 = ({(operation_194_2974[7:0])});
    assign operation_194_2945 = ({(operation_194_2973[7:0])});
    assign operation_194_2947 = ((control_194_12)?(lookup_sbox_31_output):(operation_194_2947_latch));
    assign operation_194_2948 = ((control_194_11)?(lookup_sbox_31_output):(operation_194_2948_latch));
    assign operation_194_2949 = ({(operation_194_2970[7:0])});
    assign operation_194_2950 = ({(operation_194_2965[7:0])});
    assign operation_194_2951 = ({(operation_194_2968[7:0])});
    assign operation_194_2952 = ({(operation_194_2971[7:0])});
    assign operation_194_2953 = ({(operation_194_2966[7:0])});
    assign operation_194_2954 = ({(operation_194_2969[7:0])});
    assign operation_194_2955 = ({(operation_194_2972[7:0])});
    assign operation_194_2956 = ({(operation_194_2967[7:0])});
    assign operation_194_2957 = ((control_194_20)?(lookup_sbox_31_output):(operation_194_2957_latch));
    assign operation_194_2958 = ((control_194_20)?(lookup_sbox_30_output):(operation_194_2958_latch));
    assign operation_194_2959 = ((control_194_20)?(lookup_sbox_29_output):(operation_194_2959_latch));
    assign operation_194_2960 = ((control_194_20)?(lookup_sbox_28_output):(operation_194_2960_latch));
    assign operation_194_2961 = ((control_194_20)?(lookup_sbox_27_output):(operation_194_2961_latch));
    assign operation_194_2962 = ((control_194_20)?(lookup_sbox_26_output):(operation_194_2962_latch));
    assign operation_194_2963 = ((control_194_20)?(lookup_sbox_25_output):(operation_194_2963_latch));
    assign operation_194_2964 = ((control_194_20)?(lookup_sbox_24_output):(operation_194_2964_latch));
    assign operation_194_2965 = ((control_194_20)?(lookup_sbox_23_output):(operation_194_2965_latch));
    assign operation_194_2966 = ((control_194_20)?(lookup_sbox_22_output):(operation_194_2966_latch));
    assign operation_194_2967 = ((control_194_20)?(lookup_sbox_21_output):(operation_194_2967_latch));
    assign operation_194_2968 = ((control_194_20)?(lookup_sbox_20_output):(operation_194_2968_latch));
    assign operation_194_2969 = ((control_194_20)?(lookup_sbox_19_output):(operation_194_2969_latch));
    assign operation_194_2970 = ((control_194_20)?(lookup_sbox_18_output):(operation_194_2970_latch));
    assign operation_194_2971 = ((control_194_20)?(lookup_sbox_17_output):(operation_194_2971_latch));
    assign operation_194_2972 = ((control_194_20)?(lookup_sbox_16_output):(operation_194_2972_latch));
    assign operation_194_2973 = ((control_194_11)?(lookup_sbox_30_output):(operation_194_2973_latch));
    assign operation_194_2974 = ((control_194_12)?(lookup_sbox_30_output):(operation_194_2974_latch));
    assign operation_194_2128 = (operation_194_2129);
    assign operation_194_2130 = ({(operation_194_2132[7:0])});
    assign operation_194_2132 = (operation_194_2133);
    assign operation_194_2134 = (operation_194_2135);
    assign operation_194_2136 = (operation_194_2137);
    assign operation_194_2138 = (operation_194_2139);
    assign operation_194_2140 = (operation_194_2141);
    assign operation_194_2142 = (operation_194_2143);
    assign operation_194_2144 = (operation_194_2145);
    assign operation_194_2146 = (operation_194_2147);
    assign operation_194_2148 = ({(operation_194_2226[7:0])});
    assign operation_194_2149 = ({(operation_194_2172[7:0])});
    assign operation_194_2150 = ({(operation_194_2170[7:0])});
    assign operation_194_2151 = ({(operation_194_2168[7:0])});
    assign operation_194_2152 = ({(operation_194_2166[7:0])});
    assign operation_194_2153 = ({(operation_194_2164[7:0])});
    assign operation_194_2154 = ({(operation_194_2162[7:0])});
    assign operation_194_2155 = ({(operation_194_2160[7:0])});
    assign operation_194_2156 = ({(operation_194_2158[7:0])});
    assign operation_194_2157 = ({(operation_194_2224[7:0])});
    assign operation_194_2158 = (operation_194_2159);
    assign operation_194_2160 = (operation_194_2161);
    assign operation_194_2162 = (operation_194_2163);
    assign operation_194_2164 = (operation_194_2165);
    assign operation_194_2166 = (operation_194_2167);
    assign operation_194_2168 = (operation_194_2169);
    assign operation_194_2170 = (operation_194_2171);
    assign operation_194_2172 = (operation_194_2173);
    assign operation_194_2174 = (operation_194_2175);
    assign operation_194_2176 = (operation_194_2177);
    assign operation_194_2178 = (operation_194_2179);
    assign operation_194_2180 = (operation_194_2181);
    assign operation_194_2182 = (operation_194_2183);
    assign operation_194_2184 = (operation_194_2185);
    assign operation_194_2186 = (operation_194_2187);
    assign operation_194_2188 = (operation_194_2189);
    assign operation_194_2190 = ({(operation_194_2256[7:0])});
    assign operation_194_2191 = ({(operation_194_2222[7:0])});
    assign operation_194_2192 = ({(operation_194_2254[7:0])});
    assign operation_194_2193 = ({(operation_194_2220[7:0])});
    assign operation_194_2194 = ({(operation_194_2218[7:0])});
    assign operation_194_2195 = ({(operation_194_2216[7:0])});
    assign operation_194_2196 = ({(operation_194_2214[7:0])});
    assign operation_194_2197 = ({(operation_194_2212[7:0])});
    assign operation_194_2198 = ({(operation_194_2210[7:0])});
    assign operation_194_2199 = ({(operation_194_2208[7:0])});
    assign operation_194_2200 = ({(operation_194_2252[7:0])});
    assign operation_194_2201 = ({(operation_194_2250[7:0])});
    assign operation_194_2202 = ({(operation_194_2248[7:0])});
    assign operation_194_2203 = ({(operation_194_2246[7:0])});
    assign operation_194_2204 = ({(operation_194_2244[7:0])});
    assign operation_194_2205 = ({(operation_194_2242[7:0])});
    assign operation_194_2206 = ({(operation_194_2240[7:0])});
    assign operation_194_2207 = ({(operation_194_2238[7:0])});
    assign operation_194_2208 = (operation_194_2209);
    assign operation_194_2210 = (operation_194_2211);
    assign operation_194_2212 = (operation_194_2213);
    assign operation_194_2214 = (operation_194_2215);
    assign operation_194_2216 = (operation_194_2217);
    assign operation_194_2218 = (operation_194_2219);
    assign operation_194_2220 = (operation_194_2221);
    assign operation_194_2222 = (operation_194_2223);
    assign operation_194_2224 = (operation_194_2225);
    assign operation_194_2226 = (operation_194_2227);
    assign operation_194_2228 = ({(operation_194_2286[7:0])});
    assign operation_194_2229 = ({(operation_194_2284[7:0])});
    assign operation_194_2230 = ({(operation_194_2282[7:0])});
    assign operation_194_2231 = ({(operation_194_2280[7:0])});
    assign operation_194_2232 = ({(operation_194_2278[7:0])});
    assign operation_194_2233 = ({(operation_194_2276[7:0])});
    assign operation_194_2234 = ({(operation_194_2274[7:0])});
    assign operation_194_2235 = ({(operation_194_2272[7:0])});
    assign operation_194_2236 = ({(operation_194_2270[7:0])});
    assign operation_194_2237 = ({(operation_194_2268[7:0])});
    assign operation_194_2238 = (operation_194_2239);
    assign operation_194_2240 = (operation_194_2241);
    assign operation_194_2242 = (operation_194_2243);
    assign operation_194_2244 = (operation_194_2245);
    assign operation_194_2246 = (operation_194_2247);
    assign operation_194_2248 = (operation_194_2249);
    assign operation_194_2250 = (operation_194_2251);
    assign operation_194_2252 = (operation_194_2253);
    assign operation_194_2254 = (operation_194_2255);
    assign operation_194_2256 = (operation_194_2257);
    assign operation_194_2258 = ({(operation_194_2324[7:0])});
    assign operation_194_2259 = ({(operation_194_2322[7:0])});
    assign operation_194_2260 = ({(operation_194_2319[7:0])});
    assign operation_194_2261 = ({(operation_194_2316[7:0])});
    assign operation_194_2262 = ({(operation_194_2313[7:0])});
    assign operation_194_2263 = ({(operation_194_2310[7:0])});
    assign operation_194_2264 = ({(operation_194_2307[7:0])});
    assign operation_194_2265 = ({(operation_194_2304[7:0])});
    assign operation_194_2266 = ({(operation_194_2301[7:0])});
    assign operation_194_2267 = ({(operation_194_2298[7:0])});
    assign operation_194_2268 = (operation_194_2269);
    assign operation_194_2270 = (operation_194_2271);
    assign operation_194_2272 = (operation_194_2273);
    assign operation_194_2274 = (operation_194_2275);
    assign operation_194_2276 = (operation_194_2277);
    assign operation_194_2278 = (operation_194_2279);
    assign operation_194_2280 = (operation_194_2281);
    assign operation_194_2282 = (operation_194_2283);
    assign operation_194_2284 = (operation_194_2285);
    assign operation_194_2286 = (operation_194_2287);
    assign operation_194_2288 = ({(operation_194_2386[7:0])});
    assign operation_194_2289 = ({(operation_194_2384[7:0])});
    assign operation_194_2290 = ({(operation_194_2381[7:0])});
    assign operation_194_2291 = ({(operation_194_2378[7:0])});
    assign operation_194_2292 = ({(operation_194_2375[7:0])});
    assign operation_194_2293 = ({(operation_194_2372[7:0])});
    assign operation_194_2294 = ({(operation_194_2369[7:0])});
    assign operation_194_2295 = ({(operation_194_2366[7:0])});
    assign operation_194_2296 = ({(operation_194_2363[7:0])});
    assign operation_194_2297 = ({(operation_194_2360[7:0])});
    assign operation_194_2298 = (operation_194_2299);
    assign operation_194_2301 = (operation_194_2302);
    assign operation_194_2304 = (operation_194_2305);
    assign operation_194_2307 = (operation_194_2308);
    assign operation_194_2310 = (operation_194_2311);
    assign operation_194_2313 = (operation_194_2314);
    assign operation_194_2316 = (operation_194_2317);
    assign operation_194_2319 = (operation_194_2320);
    assign operation_194_2322 = (operation_194_2323);
    assign operation_194_2324 = (operation_194_2325);
    assign operation_194_2326 = ({(operation_194_2444[7:0])});
    assign operation_194_2327 = ({(operation_194_2442[7:0])});
    assign operation_194_2331 = ({(operation_194_2434[7:0])});
    assign operation_194_2335 = ({(operation_194_2433[7:0])});
    assign operation_194_2339 = ({(operation_194_2431[7:0])});
    assign operation_194_2343 = ({(operation_194_2430[7:0])});
    assign operation_194_2347 = ({(operation_194_2428[7:0])});
    assign operation_194_2351 = ({(operation_194_2427[7:0])});
    assign operation_194_2355 = ({(operation_194_2425[7:0])});
    assign operation_194_2359 = ({(operation_194_2424[7:0])});
    assign operation_194_2360 = (operation_194_2361);
    assign operation_194_2363 = (operation_194_2364);
    assign operation_194_2366 = (operation_194_2367);
    assign operation_194_2369 = (operation_194_2370);
    assign operation_194_2372 = (operation_194_2373);
    assign operation_194_2375 = (operation_194_2376);
    assign operation_194_2378 = (operation_194_2379);
    assign operation_194_2381 = (operation_194_2382);
    assign operation_194_2384 = (operation_194_2385);
    assign operation_194_2386 = (operation_194_2387);
    assign operation_194_2388 = ({(operation_194_2475[7:0])});
    assign operation_194_2389 = ({(operation_194_2440[7:0])});
    assign operation_194_2390 = ({(operation_194_2438[7:0])});
    assign operation_194_2391 = ({(operation_194_2436[7:0])});
    assign operation_194_2395 = ({(operation_194_2469[7:0])});
    assign operation_194_2399 = ({(operation_194_2467[7:0])});
    assign operation_194_2403 = ({(operation_194_2465[7:0])});
    assign operation_194_2407 = ({(operation_194_2463[7:0])});
    assign operation_194_2411 = ({(operation_194_2461[7:0])});
    assign operation_194_2415 = ({(operation_194_2459[7:0])});
    assign operation_194_2419 = ({(operation_194_2457[7:0])});
    assign operation_194_2423 = ({(operation_194_2455[7:0])});
    assign operation_194_2424 = (operation_194_2454);
    assign operation_194_2425 = (operation_194_2426);
    assign operation_194_2427 = (operation_194_2489);
    assign operation_194_2428 = (operation_194_2429);
    assign operation_194_2430 = (operation_194_2452);
    assign operation_194_2431 = (operation_194_2432);
    assign operation_194_2433 = (operation_194_2487);
    assign operation_194_2434 = (operation_194_2435);
    assign operation_194_2436 = (operation_194_2437);
    assign operation_194_2438 = (operation_194_2439);
    assign operation_194_2440 = (operation_194_2441);
    assign operation_194_2442 = (operation_194_2443);
    assign operation_194_2444 = (operation_194_2445);
    assign operation_194_2446 = ({(operation_194_2502[7:0])});
    assign operation_194_2447 = ({(operation_194_2500[7:0])});
    assign operation_194_2448 = ({(operation_194_2519[7:0])});
    assign operation_194_2449 = ({(operation_194_2473[7:0])});
    assign operation_194_2450 = ({(operation_194_2471[7:0])});
    assign operation_194_2455 = (operation_194_2456);
    assign operation_194_2457 = (operation_194_2458);
    assign operation_194_2459 = (operation_194_2460);
    assign operation_194_2461 = (operation_194_2462);
    assign operation_194_2463 = (operation_194_2464);
    assign operation_194_2465 = (operation_194_2466);
    assign operation_194_2467 = (operation_194_2468);
    assign operation_194_2469 = (operation_194_2470);
    assign operation_194_2471 = (operation_194_2472);
    assign operation_194_2473 = (operation_194_2474);
    assign operation_194_2475 = (operation_194_2476);
    assign operation_194_2483 = ({(operation_194_2518[7:0])});
    assign operation_194_2490 = ({(operation_194_2529[7:0])});
    assign operation_194_2491 = ({(operation_194_2532[7:0])});
    assign operation_194_2492 = ({(operation_194_2531[7:0])});
    assign operation_194_2493 = ({(operation_194_2534[7:0])});
    assign operation_194_2494 = ({(operation_194_2533[7:0])});
    assign operation_194_2495 = ({(operation_194_2528[7:0])});
    assign operation_194_2496 = ({(operation_194_2535[7:0])});
    assign operation_194_2497 = ({(operation_194_2530[7:0])});
    assign operation_194_2500 = (operation_194_2501);
    assign operation_194_2502 = (operation_194_2503);
    assign operation_194_2514 = ({(operation_194_2545[7:0])});
    assign operation_194_2516 = ({(operation_194_2544[7:0])});
    assign operation_194_2518 = ((control_194_6)?(lookup_sbox_31_output):(operation_194_2518_latch));
    assign operation_194_2519 = ((control_194_6)?(lookup_sbox_30_output):(operation_194_2519_latch));
    assign operation_194_2520 = ({(operation_194_2541[7:0])});
    assign operation_194_2521 = ({(operation_194_2536[7:0])});
    assign operation_194_2522 = ({(operation_194_2539[7:0])});
    assign operation_194_2523 = ({(operation_194_2542[7:0])});
    assign operation_194_2524 = ({(operation_194_2537[7:0])});
    assign operation_194_2525 = ({(operation_194_2540[7:0])});
    assign operation_194_2526 = ({(operation_194_2543[7:0])});
    assign operation_194_2527 = ({(operation_194_2538[7:0])});
    assign operation_194_2528 = ((control_194_11)?(lookup_sbox_29_output):(operation_194_2528_latch));
    assign operation_194_2529 = ((control_194_11)?(lookup_sbox_28_output):(operation_194_2529_latch));
    assign operation_194_2530 = ((control_194_11)?(lookup_sbox_27_output):(operation_194_2530_latch));
    assign operation_194_2531 = ((control_194_11)?(lookup_sbox_26_output):(operation_194_2531_latch));
    assign operation_194_2532 = ((control_194_11)?(lookup_sbox_25_output):(operation_194_2532_latch));
    assign operation_194_2533 = ((control_194_11)?(lookup_sbox_24_output):(operation_194_2533_latch));
    assign operation_194_2534 = ((control_194_11)?(lookup_sbox_23_output):(operation_194_2534_latch));
    assign operation_194_2535 = ((control_194_11)?(lookup_sbox_22_output):(operation_194_2535_latch));
    assign operation_194_2536 = ((control_194_11)?(lookup_sbox_21_output):(operation_194_2536_latch));
    assign operation_194_2537 = ((control_194_11)?(lookup_sbox_20_output):(operation_194_2537_latch));
    assign operation_194_2538 = ((control_194_11)?(lookup_sbox_19_output):(operation_194_2538_latch));
    assign operation_194_2539 = ((control_194_11)?(lookup_sbox_18_output):(operation_194_2539_latch));
    assign operation_194_2540 = ((control_194_11)?(lookup_sbox_17_output):(operation_194_2540_latch));
    assign operation_194_2541 = ((control_194_11)?(lookup_sbox_16_output):(operation_194_2541_latch));
    assign operation_194_2542 = ((control_194_11)?(lookup_sbox_15_output):(operation_194_2542_latch));
    assign operation_194_2543 = ((control_194_11)?(lookup_sbox_14_output):(operation_194_2543_latch));
    assign operation_194_2544 = ((control_194_6)?(lookup_sbox_29_output):(operation_194_2544_latch));
    assign operation_194_2545 = ((control_194_7)?(lookup_sbox_31_output):(operation_194_2545_latch));
    assign operation_194_1699 = (operation_194_1700);
    assign operation_194_1701 = ({(operation_194_1703[7:0])});
    assign operation_194_1703 = (operation_194_1704);
    assign operation_194_1705 = (operation_194_1706);
    assign operation_194_1707 = (operation_194_1708);
    assign operation_194_1709 = (operation_194_1710);
    assign operation_194_1711 = (operation_194_1712);
    assign operation_194_1713 = (operation_194_1714);
    assign operation_194_1715 = (operation_194_1716);
    assign operation_194_1717 = (operation_194_1718);
    assign operation_194_1719 = ({(operation_194_1797[7:0])});
    assign operation_194_1720 = ({(operation_194_1743[7:0])});
    assign operation_194_1721 = ({(operation_194_1741[7:0])});
    assign operation_194_1722 = ({(operation_194_1739[7:0])});
    assign operation_194_1723 = ({(operation_194_1737[7:0])});
    assign operation_194_1724 = ({(operation_194_1735[7:0])});
    assign operation_194_1725 = ({(operation_194_1733[7:0])});
    assign operation_194_1726 = ({(operation_194_1731[7:0])});
    assign operation_194_1727 = ({(operation_194_1729[7:0])});
    assign operation_194_1728 = ({(operation_194_1795[7:0])});
    assign operation_194_1729 = (operation_194_1730);
    assign operation_194_1731 = (operation_194_1732);
    assign operation_194_1733 = (operation_194_1734);
    assign operation_194_1735 = (operation_194_1736);
    assign operation_194_1737 = (operation_194_1738);
    assign operation_194_1739 = (operation_194_1740);
    assign operation_194_1741 = (operation_194_1742);
    assign operation_194_1743 = (operation_194_1744);
    assign operation_194_1745 = (operation_194_1746);
    assign operation_194_1747 = (operation_194_1748);
    assign operation_194_1749 = (operation_194_1750);
    assign operation_194_1751 = (operation_194_1752);
    assign operation_194_1753 = (operation_194_1754);
    assign operation_194_1755 = (operation_194_1756);
    assign operation_194_1757 = (operation_194_1758);
    assign operation_194_1759 = (operation_194_1760);
    assign operation_194_1761 = ({(operation_194_1827[7:0])});
    assign operation_194_1762 = ({(operation_194_1793[7:0])});
    assign operation_194_1763 = ({(operation_194_1825[7:0])});
    assign operation_194_1764 = ({(operation_194_1791[7:0])});
    assign operation_194_1765 = ({(operation_194_1789[7:0])});
    assign operation_194_1766 = ({(operation_194_1787[7:0])});
    assign operation_194_1767 = ({(operation_194_1785[7:0])});
    assign operation_194_1768 = ({(operation_194_1783[7:0])});
    assign operation_194_1769 = ({(operation_194_1781[7:0])});
    assign operation_194_1770 = ({(operation_194_1779[7:0])});
    assign operation_194_1771 = ({(operation_194_1823[7:0])});
    assign operation_194_1772 = ({(operation_194_1821[7:0])});
    assign operation_194_1773 = ({(operation_194_1819[7:0])});
    assign operation_194_1774 = ({(operation_194_1817[7:0])});
    assign operation_194_1775 = ({(operation_194_1815[7:0])});
    assign operation_194_1776 = ({(operation_194_1813[7:0])});
    assign operation_194_1777 = ({(operation_194_1811[7:0])});
    assign operation_194_1778 = ({(operation_194_1809[7:0])});
    assign operation_194_1779 = (operation_194_1780);
    assign operation_194_1781 = (operation_194_1782);
    assign operation_194_1783 = (operation_194_1784);
    assign operation_194_1785 = (operation_194_1786);
    assign operation_194_1787 = (operation_194_1788);
    assign operation_194_1789 = (operation_194_1790);
    assign operation_194_1791 = (operation_194_1792);
    assign operation_194_1793 = (operation_194_1794);
    assign operation_194_1795 = (operation_194_1796);
    assign operation_194_1797 = (operation_194_1798);
    assign operation_194_1799 = ({(operation_194_1857[7:0])});
    assign operation_194_1800 = ({(operation_194_1855[7:0])});
    assign operation_194_1801 = ({(operation_194_1853[7:0])});
    assign operation_194_1802 = ({(operation_194_1851[7:0])});
    assign operation_194_1803 = ({(operation_194_1849[7:0])});
    assign operation_194_1804 = ({(operation_194_1847[7:0])});
    assign operation_194_1805 = ({(operation_194_1845[7:0])});
    assign operation_194_1806 = ({(operation_194_1843[7:0])});
    assign operation_194_1807 = ({(operation_194_1841[7:0])});
    assign operation_194_1808 = ({(operation_194_1839[7:0])});
    assign operation_194_1809 = (operation_194_1810);
    assign operation_194_1811 = (operation_194_1812);
    assign operation_194_1813 = (operation_194_1814);
    assign operation_194_1815 = (operation_194_1816);
    assign operation_194_1817 = (operation_194_1818);
    assign operation_194_1819 = (operation_194_1820);
    assign operation_194_1821 = (operation_194_1822);
    assign operation_194_1823 = (operation_194_1824);
    assign operation_194_1825 = (operation_194_1826);
    assign operation_194_1827 = (operation_194_1828);
    assign operation_194_1829 = ({(operation_194_1895[7:0])});
    assign operation_194_1830 = ({(operation_194_1893[7:0])});
    assign operation_194_1831 = ({(operation_194_1890[7:0])});
    assign operation_194_1832 = ({(operation_194_1887[7:0])});
    assign operation_194_1833 = ({(operation_194_1884[7:0])});
    assign operation_194_1834 = ({(operation_194_1881[7:0])});
    assign operation_194_1835 = ({(operation_194_1878[7:0])});
    assign operation_194_1836 = ({(operation_194_1875[7:0])});
    assign operation_194_1837 = ({(operation_194_1872[7:0])});
    assign operation_194_1838 = ({(operation_194_1869[7:0])});
    assign operation_194_1839 = (operation_194_1840);
    assign operation_194_1841 = (operation_194_1842);
    assign operation_194_1843 = (operation_194_1844);
    assign operation_194_1845 = (operation_194_1846);
    assign operation_194_1847 = (operation_194_1848);
    assign operation_194_1849 = (operation_194_1850);
    assign operation_194_1851 = (operation_194_1852);
    assign operation_194_1853 = (operation_194_1854);
    assign operation_194_1855 = (operation_194_1856);
    assign operation_194_1857 = (operation_194_1858);
    assign operation_194_1859 = ({(operation_194_1957[7:0])});
    assign operation_194_1860 = ({(operation_194_1955[7:0])});
    assign operation_194_1861 = ({(operation_194_1952[7:0])});
    assign operation_194_1862 = ({(operation_194_1949[7:0])});
    assign operation_194_1863 = ({(operation_194_1946[7:0])});
    assign operation_194_1864 = ({(operation_194_1943[7:0])});
    assign operation_194_1865 = ({(operation_194_1940[7:0])});
    assign operation_194_1866 = ({(operation_194_1937[7:0])});
    assign operation_194_1867 = ({(operation_194_1934[7:0])});
    assign operation_194_1868 = ({(operation_194_1931[7:0])});
    assign operation_194_1869 = (operation_194_1870);
    assign operation_194_1872 = (operation_194_1873);
    assign operation_194_1875 = (operation_194_1876);
    assign operation_194_1878 = (operation_194_1879);
    assign operation_194_1881 = (operation_194_1882);
    assign operation_194_1884 = (operation_194_1885);
    assign operation_194_1887 = (operation_194_1888);
    assign operation_194_1890 = (operation_194_1891);
    assign operation_194_1893 = (operation_194_1894);
    assign operation_194_1895 = (operation_194_1896);
    assign operation_194_1897 = ({(operation_194_2015[7:0])});
    assign operation_194_1898 = ({(operation_194_2013[7:0])});
    assign operation_194_1902 = ({(operation_194_2005[7:0])});
    assign operation_194_1906 = ({(operation_194_2004[7:0])});
    assign operation_194_1910 = ({(operation_194_2002[7:0])});
    assign operation_194_1914 = ({(operation_194_2001[7:0])});
    assign operation_194_1918 = ({(operation_194_1999[7:0])});
    assign operation_194_1922 = ({(operation_194_1998[7:0])});
    assign operation_194_1926 = ({(operation_194_1996[7:0])});
    assign operation_194_1930 = ({(operation_194_1995[7:0])});
    assign operation_194_1931 = (operation_194_1932);
    assign operation_194_1934 = (operation_194_1935);
    assign operation_194_1937 = (operation_194_1938);
    assign operation_194_1940 = (operation_194_1941);
    assign operation_194_1943 = (operation_194_1944);
    assign operation_194_1946 = (operation_194_1947);
    assign operation_194_1949 = (operation_194_1950);
    assign operation_194_1952 = (operation_194_1953);
    assign operation_194_1955 = (operation_194_1956);
    assign operation_194_1957 = (operation_194_1958);
    assign operation_194_1959 = ({(operation_194_2046[7:0])});
    assign operation_194_1960 = ({(operation_194_2011[7:0])});
    assign operation_194_1961 = ({(operation_194_2009[7:0])});
    assign operation_194_1962 = ({(operation_194_2007[7:0])});
    assign operation_194_1966 = ({(operation_194_2040[7:0])});
    assign operation_194_1970 = ({(operation_194_2038[7:0])});
    assign operation_194_1974 = ({(operation_194_2036[7:0])});
    assign operation_194_1978 = ({(operation_194_2034[7:0])});
    assign operation_194_1982 = ({(operation_194_2032[7:0])});
    assign operation_194_1986 = ({(operation_194_2030[7:0])});
    assign operation_194_1990 = ({(operation_194_2028[7:0])});
    assign operation_194_1994 = ({(operation_194_2026[7:0])});
    assign operation_194_1995 = (operation_194_2025);
    assign operation_194_1996 = (operation_194_1997);
    assign operation_194_1998 = (operation_194_2060);
    assign operation_194_1999 = (operation_194_2000);
    assign operation_194_2001 = (operation_194_2023);
    assign operation_194_2002 = (operation_194_2003);
    assign operation_194_2004 = (operation_194_2058);
    assign operation_194_2005 = (operation_194_2006);
    assign operation_194_2007 = (operation_194_2008);
    assign operation_194_2009 = (operation_194_2010);
    assign operation_194_2011 = (operation_194_2012);
    assign operation_194_2013 = (operation_194_2014);
    assign operation_194_2015 = (operation_194_2016);
    assign operation_194_2017 = ({(operation_194_2073[7:0])});
    assign operation_194_2018 = ({(operation_194_2071[7:0])});
    assign operation_194_2019 = ({(operation_194_2090[7:0])});
    assign operation_194_2020 = ({(operation_194_2044[7:0])});
    assign operation_194_2021 = ({(operation_194_2042[7:0])});
    assign operation_194_2026 = (operation_194_2027);
    assign operation_194_2028 = (operation_194_2029);
    assign operation_194_2030 = (operation_194_2031);
    assign operation_194_2032 = (operation_194_2033);
    assign operation_194_2034 = (operation_194_2035);
    assign operation_194_2036 = (operation_194_2037);
    assign operation_194_2038 = (operation_194_2039);
    assign operation_194_2040 = (operation_194_2041);
    assign operation_194_2042 = (operation_194_2043);
    assign operation_194_2044 = (operation_194_2045);
    assign operation_194_2046 = (operation_194_2047);
    assign operation_194_2054 = ({(operation_194_2089[7:0])});
    assign operation_194_2061 = ({(operation_194_2100[7:0])});
    assign operation_194_2062 = ({(operation_194_2103[7:0])});
    assign operation_194_2063 = ({(operation_194_2102[7:0])});
    assign operation_194_2064 = ({(operation_194_2105[7:0])});
    assign operation_194_2065 = ({(operation_194_2104[7:0])});
    assign operation_194_2066 = ({(operation_194_2099[7:0])});
    assign operation_194_2067 = ({(operation_194_2106[7:0])});
    assign operation_194_2068 = ({(operation_194_2101[7:0])});
    assign operation_194_2071 = (operation_194_2072);
    assign operation_194_2073 = (operation_194_2074);
    assign operation_194_2085 = ({(operation_194_2116[7:0])});
    assign operation_194_2087 = ({(operation_194_2115[7:0])});
    assign operation_194_2089 = ((control_194_1)?(lookup_sbox_31_output):(operation_194_2089_latch));
    assign operation_194_2090 = ((control_194_1)?(lookup_sbox_30_output):(operation_194_2090_latch));
    assign operation_194_2091 = ({(operation_194_2112[7:0])});
    assign operation_194_2092 = ({(operation_194_2107[7:0])});
    assign operation_194_2093 = ({(operation_194_2110[7:0])});
    assign operation_194_2094 = ({(operation_194_2113[7:0])});
    assign operation_194_2095 = ({(operation_194_2108[7:0])});
    assign operation_194_2096 = ({(operation_194_2111[7:0])});
    assign operation_194_2097 = ({(operation_194_2114[7:0])});
    assign operation_194_2098 = ({(operation_194_2109[7:0])});
    assign operation_194_2099 = ((control_194_2)?(lookup_sbox_31_output):(operation_194_2099_latch));
    assign operation_194_2100 = ((control_194_2)?(lookup_sbox_30_output):(operation_194_2100_latch));
    assign operation_194_2101 = ((control_194_2)?(lookup_sbox_29_output):(operation_194_2101_latch));
    assign operation_194_2102 = ((control_194_2)?(lookup_sbox_28_output):(operation_194_2102_latch));
    assign operation_194_2103 = ((control_194_2)?(lookup_sbox_27_output):(operation_194_2103_latch));
    assign operation_194_2104 = ((control_194_2)?(lookup_sbox_26_output):(operation_194_2104_latch));
    assign operation_194_2105 = ((control_194_2)?(lookup_sbox_25_output):(operation_194_2105_latch));
    assign operation_194_2106 = ((control_194_2)?(lookup_sbox_24_output):(operation_194_2106_latch));
    assign operation_194_2107 = ((control_194_2)?(lookup_sbox_23_output):(operation_194_2107_latch));
    assign operation_194_2108 = ((control_194_2)?(lookup_sbox_22_output):(operation_194_2108_latch));
    assign operation_194_2109 = ((control_194_2)?(lookup_sbox_21_output):(operation_194_2109_latch));
    assign operation_194_2110 = ((control_194_2)?(lookup_sbox_20_output):(operation_194_2110_latch));
    assign operation_194_2111 = ((control_194_2)?(lookup_sbox_19_output):(operation_194_2111_latch));
    assign operation_194_2112 = ((control_194_2)?(lookup_sbox_18_output):(operation_194_2112_latch));
    assign operation_194_2113 = ((control_194_2)?(lookup_sbox_17_output):(operation_194_2113_latch));
    assign operation_194_2114 = ((control_194_2)?(lookup_sbox_16_output):(operation_194_2114_latch));
    assign operation_194_2115 = ((control_194_1)?(lookup_sbox_29_output):(operation_194_2115_latch));
    assign operation_194_2116 = ((control_194_1)?(lookup_sbox_28_output):(operation_194_2116_latch));
    assign operation_194_127 = (operation_194_126);
    assign operation_194_123 = ({(operation_194_122[127:120])});
    assign operation_194_7 = (operation_194_6);
    assign operation_194_23 = (operation_194_22);
    assign operation_194_39 = (operation_194_38);
    assign operation_194_55 = (operation_194_54);
    assign operation_194_71 = (operation_194_70);
    assign operation_194_87 = (operation_194_86);
    assign operation_194_103 = (operation_194_102);
    assign operation_194_119 = (operation_194_118);
    assign operation_194_117 = ({(operation_194_124[119:112])});
    assign operation_194_115 = ({(operation_194_122[119:112])});
    assign operation_194_101 = ({(operation_194_124[103:96])});
    assign operation_194_99 = ({(operation_194_122[103:96])});
    assign operation_194_85 = ({(operation_194_124[87:80])});
    assign operation_194_83 = ({(operation_194_122[87:80])});
    assign operation_194_69 = ({(operation_194_124[71:64])});
    assign operation_194_67 = ({(operation_194_122[71:64])});
    assign operation_194_53 = ({(operation_194_124[55:48])});
    assign operation_194_51 = ({(operation_194_122[55:48])});
    assign operation_194_37 = ({(operation_194_124[39:32])});
    assign operation_194_35 = ({(operation_194_122[39:32])});
    assign operation_194_21 = ({(operation_194_124[23:16])});
    assign operation_194_19 = ({(operation_194_122[23:16])});
    assign operation_194_5 = ({(operation_194_124[7:0])});
    assign operation_194_3 = ({(operation_194_122[7:0])});
    assign operation_194_15 = (operation_194_14);
    assign operation_194_11 = ({(operation_194_122[15:8])});
    assign operation_194_13 = ({(operation_194_124[15:8])});
    assign operation_194_31 = (operation_194_30);
    assign operation_194_27 = ({(operation_194_122[31:24])});
    assign operation_194_29 = ({(operation_194_124[31:24])});
    assign operation_194_47 = (operation_194_46);
    assign operation_194_43 = ({(operation_194_122[47:40])});
    assign operation_194_45 = ({(operation_194_124[47:40])});
    assign operation_194_63 = (operation_194_62);
    assign operation_194_59 = ({(operation_194_122[63:56])});
    assign operation_194_61 = ({(operation_194_124[63:56])});
    assign operation_194_79 = (operation_194_78);
    assign operation_194_75 = ({(operation_194_122[79:72])});
    assign operation_194_77 = ({(operation_194_124[79:72])});
    assign operation_194_95 = (operation_194_94);
    assign operation_194_91 = ({(operation_194_122[95:88])});
    assign operation_194_93 = ({(operation_194_124[95:88])});
    assign operation_194_111 = (operation_194_110);
    assign operation_194_107 = ({(operation_194_122[111:104])});
    assign operation_194_109 = ({(operation_194_124[111:104])});
    assign operation_194_125 = ({(operation_194_124[127:120])});
    assign operation_194_5601 = (32'd54);
    assign operation_194_5597 = (32'd27);
    assign operation_194_5592 = (32'd128);
    assign operation_194_5587 = (32'd64);
    assign operation_194_5582 = (32'd32);
    assign operation_194_5577 = (32'd16);
    assign operation_194_5572 = (32'd8);
    assign operation_194_5567 = (32'd4);
    assign operation_194_5562 = (32'd2);
    assign operation_194_5557 = (32'd1);
    assign operation_194_2119 = (32'd7);
    assign operation_194_124 = (input_key_194);
    assign operation_194_122 = (input_in_194);
    assign control_194_end = (control_194_83);
    assign control_194_0 = (control_194_start);
    
    always_ff @(posedge clk)
    if(rst)
         begin
            finish <= 1'd0;
            AES128_encrypt <= 128'd0;
            operation_194_1664 <= 32'd0;
            operation_194_1536 <= 32'd0;
            operation_194_1680 <= 32'd0;
            operation_194_1632 <= 32'd0;
            operation_194_1672 <= 32'd0;
            operation_194_1688 <= 32'd0;
            operation_194_1504 <= 32'd0;
            operation_194_1552 <= 32'd0;
            operation_194_1648 <= 32'd0;
            operation_194_1600 <= 32'd0;
            operation_194_1544 <= 32'd0;
            operation_194_1560 <= 32'd0;
            operation_194_1656 <= 32'd0;
            operation_194_1640 <= 32'd0;
            operation_194_1472 <= 32'd0;
            operation_194_1520 <= 32'd0;
            operation_194_1616 <= 32'd0;
            operation_194_1568 <= 32'd0;
            operation_194_1512 <= 32'd0;
            operation_194_1528 <= 32'd0;
            operation_194_1624 <= 32'd0;
            operation_194_1608 <= 32'd0;
            operation_194_1440 <= 32'd0;
            operation_194_1488 <= 32'd0;
            operation_194_1584 <= 32'd0;
            operation_194_1432 <= 32'd0;
            operation_194_1480 <= 32'd0;
            operation_194_1496 <= 32'd0;
            operation_194_1592 <= 32'd0;
            operation_194_1576 <= 32'd0;
            operation_194_1456 <= 32'd0;
            operation_194_1448 <= 32'd0;
            operation_194_1464 <= 32'd0;
            operation_194_1338_latch <= 8'd0;
            operation_194_1328_latch <= 8'd0;
            operation_194_1318_latch <= 8'd0;
            operation_194_1308_latch <= 8'd0;
            operation_194_1298_latch <= 8'd0;
            operation_194_1288_latch <= 8'd0;
            operation_194_1278_latch <= 8'd0;
            operation_194_1268_latch <= 8'd0;
            operation_194_1273_latch <= 8'd0;
            operation_194_1283_latch <= 8'd0;
            operation_194_1293_latch <= 8'd0;
            operation_194_1303_latch <= 8'd0;
            operation_194_1313_latch <= 8'd0;
            operation_194_1323_latch <= 8'd0;
            operation_194_1333_latch <= 8'd0;
            operation_194_1343_latch <= 8'd0;
            operation_194_1413_latch <= 8'd0;
            operation_194_1423_latch <= 8'd0;
            operation_194_1408_latch <= 8'd0;
            operation_194_1418_latch <= 8'd0;
            operation_194_5132 <= 32'd0;
            operation_194_5136 <= 32'd0;
            operation_194_5138 <= 32'd0;
            operation_194_5140 <= 32'd0;
            operation_194_5142 <= 32'd0;
            operation_194_5144 <= 32'd0;
            operation_194_5146 <= 32'd0;
            operation_194_5148 <= 32'd0;
            operation_194_5150 <= 32'd0;
            operation_194_5162 <= 32'd0;
            operation_194_5164 <= 32'd0;
            operation_194_5166 <= 32'd0;
            operation_194_5168 <= 32'd0;
            operation_194_5170 <= 32'd0;
            operation_194_5172 <= 32'd0;
            operation_194_5174 <= 32'd0;
            operation_194_5176 <= 32'd0;
            operation_194_5178 <= 32'd0;
            operation_194_5180 <= 32'd0;
            operation_194_5182 <= 32'd0;
            operation_194_5184 <= 32'd0;
            operation_194_5186 <= 32'd0;
            operation_194_5188 <= 32'd0;
            operation_194_5190 <= 32'd0;
            operation_194_5192 <= 32'd0;
            operation_194_5212 <= 32'd0;
            operation_194_5214 <= 32'd0;
            operation_194_5216 <= 32'd0;
            operation_194_5218 <= 32'd0;
            operation_194_5220 <= 32'd0;
            operation_194_5222 <= 32'd0;
            operation_194_5224 <= 32'd0;
            operation_194_5226 <= 32'd0;
            operation_194_5228 <= 32'd0;
            operation_194_5230 <= 32'd0;
            operation_194_5242 <= 32'd0;
            operation_194_5244 <= 32'd0;
            operation_194_5246 <= 32'd0;
            operation_194_5248 <= 32'd0;
            operation_194_5250 <= 32'd0;
            operation_194_5252 <= 32'd0;
            operation_194_5254 <= 32'd0;
            operation_194_5256 <= 32'd0;
            operation_194_5258 <= 32'd0;
            operation_194_5260 <= 32'd0;
            operation_194_5272 <= 32'd0;
            operation_194_5274 <= 32'd0;
            operation_194_5276 <= 32'd0;
            operation_194_5278 <= 32'd0;
            operation_194_5280 <= 32'd0;
            operation_194_5282 <= 32'd0;
            operation_194_5284 <= 32'd0;
            operation_194_5286 <= 32'd0;
            operation_194_5288 <= 32'd0;
            operation_194_5290 <= 32'd0;
            operation_194_5302 <= 32'd0;
            operation_194_5303 <= 32'd0;
            operation_194_5305 <= 32'd0;
            operation_194_5306 <= 32'd0;
            operation_194_5308 <= 32'd0;
            operation_194_5309 <= 32'd0;
            operation_194_5311 <= 32'd0;
            operation_194_5312 <= 32'd0;
            operation_194_5314 <= 32'd0;
            operation_194_5315 <= 32'd0;
            operation_194_5317 <= 32'd0;
            operation_194_5318 <= 32'd0;
            operation_194_5320 <= 32'd0;
            operation_194_5321 <= 32'd0;
            operation_194_5323 <= 32'd0;
            operation_194_5324 <= 32'd0;
            operation_194_5326 <= 32'd0;
            operation_194_5328 <= 32'd0;
            operation_194_5331 <= 32'd0;
            operation_194_5332 <= 32'd0;
            operation_194_5333 <= 32'd0;
            operation_194_5335 <= 32'd0;
            operation_194_5336 <= 32'd0;
            operation_194_5337 <= 32'd0;
            operation_194_5339 <= 32'd0;
            operation_194_5340 <= 32'd0;
            operation_194_5341 <= 32'd0;
            operation_194_5343 <= 32'd0;
            operation_194_5344 <= 32'd0;
            operation_194_5345 <= 32'd0;
            operation_194_5347 <= 32'd0;
            operation_194_5348 <= 32'd0;
            operation_194_5349 <= 32'd0;
            operation_194_5351 <= 32'd0;
            operation_194_5352 <= 32'd0;
            operation_194_5353 <= 32'd0;
            operation_194_5355 <= 32'd0;
            operation_194_5356 <= 32'd0;
            operation_194_5357 <= 32'd0;
            operation_194_5359 <= 32'd0;
            operation_194_5360 <= 32'd0;
            operation_194_5361 <= 32'd0;
            operation_194_5364 <= 32'd0;
            operation_194_5365 <= 32'd0;
            operation_194_5367 <= 32'd0;
            operation_194_5368 <= 32'd0;
            operation_194_5370 <= 32'd0;
            operation_194_5371 <= 32'd0;
            operation_194_5373 <= 32'd0;
            operation_194_5374 <= 32'd0;
            operation_194_5376 <= 32'd0;
            operation_194_5377 <= 32'd0;
            operation_194_5379 <= 32'd0;
            operation_194_5380 <= 32'd0;
            operation_194_5382 <= 32'd0;
            operation_194_5383 <= 32'd0;
            operation_194_5385 <= 32'd0;
            operation_194_5386 <= 32'd0;
            operation_194_5388 <= 32'd0;
            operation_194_5390 <= 32'd0;
            operation_194_5395 <= 32'd0;
            operation_194_5396 <= 32'd0;
            operation_194_5397 <= 32'd0;
            operation_194_5399 <= 32'd0;
            operation_194_5400 <= 32'd0;
            operation_194_5401 <= 32'd0;
            operation_194_5403 <= 32'd0;
            operation_194_5404 <= 32'd0;
            operation_194_5405 <= 32'd0;
            operation_194_5407 <= 32'd0;
            operation_194_5408 <= 32'd0;
            operation_194_5409 <= 32'd0;
            operation_194_5411 <= 32'd0;
            operation_194_5412 <= 32'd0;
            operation_194_5413 <= 32'd0;
            operation_194_5415 <= 32'd0;
            operation_194_5416 <= 32'd0;
            operation_194_5417 <= 32'd0;
            operation_194_5419 <= 32'd0;
            operation_194_5420 <= 32'd0;
            operation_194_5421 <= 32'd0;
            operation_194_5423 <= 32'd0;
            operation_194_5424 <= 32'd0;
            operation_194_5425 <= 32'd0;
            operation_194_5429 <= 32'd0;
            operation_194_5432 <= 32'd0;
            operation_194_5435 <= 32'd0;
            operation_194_5438 <= 32'd0;
            operation_194_5440 <= 32'd0;
            operation_194_5442 <= 32'd0;
            operation_194_5444 <= 32'd0;
            operation_194_5446 <= 32'd0;
            operation_194_5448 <= 32'd0;
            operation_194_5454 <= 32'd0;
            operation_194_5455 <= 32'd0;
            operation_194_5456 <= 32'd0;
            operation_194_5457 <= 32'd0;
            operation_194_5459 <= 32'd0;
            operation_194_5461 <= 32'd0;
            operation_194_5463 <= 32'd0;
            operation_194_5465 <= 32'd0;
            operation_194_5467 <= 32'd0;
            operation_194_5469 <= 32'd0;
            operation_194_5471 <= 32'd0;
            operation_194_5473 <= 32'd0;
            operation_194_5475 <= 32'd0;
            operation_194_5477 <= 32'd0;
            operation_194_5479 <= 32'd0;
            operation_194_5489 <= 32'd0;
            operation_194_5490 <= 32'd0;
            operation_194_5491 <= 32'd0;
            operation_194_5492 <= 32'd0;
            operation_194_5504 <= 32'd0;
            operation_194_5506 <= 32'd0;
            operation_194_5521_latch <= 8'd0;
            operation_194_5522_latch <= 8'd0;
            operation_194_5531_latch <= 8'd0;
            operation_194_5532_latch <= 8'd0;
            operation_194_5533_latch <= 8'd0;
            operation_194_5534_latch <= 8'd0;
            operation_194_5535_latch <= 8'd0;
            operation_194_5536_latch <= 8'd0;
            operation_194_5537_latch <= 8'd0;
            operation_194_5538_latch <= 8'd0;
            operation_194_5539_latch <= 8'd0;
            operation_194_5540_latch <= 8'd0;
            operation_194_5541_latch <= 8'd0;
            operation_194_5542_latch <= 8'd0;
            operation_194_5543_latch <= 8'd0;
            operation_194_5544_latch <= 8'd0;
            operation_194_5545_latch <= 8'd0;
            operation_194_5546_latch <= 8'd0;
            operation_194_5547_latch <= 8'd0;
            operation_194_5548_latch <= 8'd0;
            operation_194_4703 <= 32'd0;
            operation_194_4707 <= 32'd0;
            operation_194_4709 <= 32'd0;
            operation_194_4711 <= 32'd0;
            operation_194_4713 <= 32'd0;
            operation_194_4715 <= 32'd0;
            operation_194_4717 <= 32'd0;
            operation_194_4719 <= 32'd0;
            operation_194_4721 <= 32'd0;
            operation_194_4733 <= 32'd0;
            operation_194_4735 <= 32'd0;
            operation_194_4737 <= 32'd0;
            operation_194_4739 <= 32'd0;
            operation_194_4741 <= 32'd0;
            operation_194_4743 <= 32'd0;
            operation_194_4745 <= 32'd0;
            operation_194_4747 <= 32'd0;
            operation_194_4749 <= 32'd0;
            operation_194_4751 <= 32'd0;
            operation_194_4753 <= 32'd0;
            operation_194_4755 <= 32'd0;
            operation_194_4757 <= 32'd0;
            operation_194_4759 <= 32'd0;
            operation_194_4761 <= 32'd0;
            operation_194_4763 <= 32'd0;
            operation_194_4783 <= 32'd0;
            operation_194_4785 <= 32'd0;
            operation_194_4787 <= 32'd0;
            operation_194_4789 <= 32'd0;
            operation_194_4791 <= 32'd0;
            operation_194_4793 <= 32'd0;
            operation_194_4795 <= 32'd0;
            operation_194_4797 <= 32'd0;
            operation_194_4799 <= 32'd0;
            operation_194_4801 <= 32'd0;
            operation_194_4813 <= 32'd0;
            operation_194_4815 <= 32'd0;
            operation_194_4817 <= 32'd0;
            operation_194_4819 <= 32'd0;
            operation_194_4821 <= 32'd0;
            operation_194_4823 <= 32'd0;
            operation_194_4825 <= 32'd0;
            operation_194_4827 <= 32'd0;
            operation_194_4829 <= 32'd0;
            operation_194_4831 <= 32'd0;
            operation_194_4843 <= 32'd0;
            operation_194_4845 <= 32'd0;
            operation_194_4847 <= 32'd0;
            operation_194_4849 <= 32'd0;
            operation_194_4851 <= 32'd0;
            operation_194_4853 <= 32'd0;
            operation_194_4855 <= 32'd0;
            operation_194_4857 <= 32'd0;
            operation_194_4859 <= 32'd0;
            operation_194_4861 <= 32'd0;
            operation_194_4873 <= 32'd0;
            operation_194_4874 <= 32'd0;
            operation_194_4876 <= 32'd0;
            operation_194_4877 <= 32'd0;
            operation_194_4879 <= 32'd0;
            operation_194_4880 <= 32'd0;
            operation_194_4882 <= 32'd0;
            operation_194_4883 <= 32'd0;
            operation_194_4885 <= 32'd0;
            operation_194_4886 <= 32'd0;
            operation_194_4888 <= 32'd0;
            operation_194_4889 <= 32'd0;
            operation_194_4891 <= 32'd0;
            operation_194_4892 <= 32'd0;
            operation_194_4894 <= 32'd0;
            operation_194_4895 <= 32'd0;
            operation_194_4897 <= 32'd0;
            operation_194_4899 <= 32'd0;
            operation_194_4902 <= 32'd0;
            operation_194_4903 <= 32'd0;
            operation_194_4904 <= 32'd0;
            operation_194_4906 <= 32'd0;
            operation_194_4907 <= 32'd0;
            operation_194_4908 <= 32'd0;
            operation_194_4910 <= 32'd0;
            operation_194_4911 <= 32'd0;
            operation_194_4912 <= 32'd0;
            operation_194_4914 <= 32'd0;
            operation_194_4915 <= 32'd0;
            operation_194_4916 <= 32'd0;
            operation_194_4918 <= 32'd0;
            operation_194_4919 <= 32'd0;
            operation_194_4920 <= 32'd0;
            operation_194_4922 <= 32'd0;
            operation_194_4923 <= 32'd0;
            operation_194_4924 <= 32'd0;
            operation_194_4926 <= 32'd0;
            operation_194_4927 <= 32'd0;
            operation_194_4928 <= 32'd0;
            operation_194_4930 <= 32'd0;
            operation_194_4931 <= 32'd0;
            operation_194_4932 <= 32'd0;
            operation_194_4935 <= 32'd0;
            operation_194_4936 <= 32'd0;
            operation_194_4938 <= 32'd0;
            operation_194_4939 <= 32'd0;
            operation_194_4941 <= 32'd0;
            operation_194_4942 <= 32'd0;
            operation_194_4944 <= 32'd0;
            operation_194_4945 <= 32'd0;
            operation_194_4947 <= 32'd0;
            operation_194_4948 <= 32'd0;
            operation_194_4950 <= 32'd0;
            operation_194_4951 <= 32'd0;
            operation_194_4953 <= 32'd0;
            operation_194_4954 <= 32'd0;
            operation_194_4956 <= 32'd0;
            operation_194_4957 <= 32'd0;
            operation_194_4959 <= 32'd0;
            operation_194_4961 <= 32'd0;
            operation_194_4966 <= 32'd0;
            operation_194_4967 <= 32'd0;
            operation_194_4968 <= 32'd0;
            operation_194_4970 <= 32'd0;
            operation_194_4971 <= 32'd0;
            operation_194_4972 <= 32'd0;
            operation_194_4974 <= 32'd0;
            operation_194_4975 <= 32'd0;
            operation_194_4976 <= 32'd0;
            operation_194_4978 <= 32'd0;
            operation_194_4979 <= 32'd0;
            operation_194_4980 <= 32'd0;
            operation_194_4982 <= 32'd0;
            operation_194_4983 <= 32'd0;
            operation_194_4984 <= 32'd0;
            operation_194_4986 <= 32'd0;
            operation_194_4987 <= 32'd0;
            operation_194_4988 <= 32'd0;
            operation_194_4990 <= 32'd0;
            operation_194_4991 <= 32'd0;
            operation_194_4992 <= 32'd0;
            operation_194_4994 <= 32'd0;
            operation_194_4995 <= 32'd0;
            operation_194_4996 <= 32'd0;
            operation_194_5000 <= 32'd0;
            operation_194_5003 <= 32'd0;
            operation_194_5006 <= 32'd0;
            operation_194_5009 <= 32'd0;
            operation_194_5011 <= 32'd0;
            operation_194_5013 <= 32'd0;
            operation_194_5015 <= 32'd0;
            operation_194_5017 <= 32'd0;
            operation_194_5019 <= 32'd0;
            operation_194_5025 <= 32'd0;
            operation_194_5026 <= 32'd0;
            operation_194_5027 <= 32'd0;
            operation_194_5028 <= 32'd0;
            operation_194_5030 <= 32'd0;
            operation_194_5032 <= 32'd0;
            operation_194_5034 <= 32'd0;
            operation_194_5036 <= 32'd0;
            operation_194_5038 <= 32'd0;
            operation_194_5040 <= 32'd0;
            operation_194_5042 <= 32'd0;
            operation_194_5044 <= 32'd0;
            operation_194_5046 <= 32'd0;
            operation_194_5048 <= 32'd0;
            operation_194_5050 <= 32'd0;
            operation_194_5060 <= 32'd0;
            operation_194_5061 <= 32'd0;
            operation_194_5062 <= 32'd0;
            operation_194_5063 <= 32'd0;
            operation_194_5075 <= 32'd0;
            operation_194_5077 <= 32'd0;
            operation_194_5092_latch <= 8'd0;
            operation_194_5093_latch <= 8'd0;
            operation_194_5102_latch <= 8'd0;
            operation_194_5103_latch <= 8'd0;
            operation_194_5104_latch <= 8'd0;
            operation_194_5105_latch <= 8'd0;
            operation_194_5106_latch <= 8'd0;
            operation_194_5107_latch <= 8'd0;
            operation_194_5108_latch <= 8'd0;
            operation_194_5109_latch <= 8'd0;
            operation_194_5110_latch <= 8'd0;
            operation_194_5111_latch <= 8'd0;
            operation_194_5112_latch <= 8'd0;
            operation_194_5113_latch <= 8'd0;
            operation_194_5114_latch <= 8'd0;
            operation_194_5115_latch <= 8'd0;
            operation_194_5116_latch <= 8'd0;
            operation_194_5117_latch <= 8'd0;
            operation_194_5118_latch <= 8'd0;
            operation_194_5119_latch <= 8'd0;
            operation_194_4274 <= 32'd0;
            operation_194_4278 <= 32'd0;
            operation_194_4280 <= 32'd0;
            operation_194_4282 <= 32'd0;
            operation_194_4284 <= 32'd0;
            operation_194_4286 <= 32'd0;
            operation_194_4288 <= 32'd0;
            operation_194_4290 <= 32'd0;
            operation_194_4292 <= 32'd0;
            operation_194_4304 <= 32'd0;
            operation_194_4306 <= 32'd0;
            operation_194_4308 <= 32'd0;
            operation_194_4310 <= 32'd0;
            operation_194_4312 <= 32'd0;
            operation_194_4314 <= 32'd0;
            operation_194_4316 <= 32'd0;
            operation_194_4318 <= 32'd0;
            operation_194_4320 <= 32'd0;
            operation_194_4322 <= 32'd0;
            operation_194_4324 <= 32'd0;
            operation_194_4326 <= 32'd0;
            operation_194_4328 <= 32'd0;
            operation_194_4330 <= 32'd0;
            operation_194_4332 <= 32'd0;
            operation_194_4334 <= 32'd0;
            operation_194_4354 <= 32'd0;
            operation_194_4356 <= 32'd0;
            operation_194_4358 <= 32'd0;
            operation_194_4360 <= 32'd0;
            operation_194_4362 <= 32'd0;
            operation_194_4364 <= 32'd0;
            operation_194_4366 <= 32'd0;
            operation_194_4368 <= 32'd0;
            operation_194_4370 <= 32'd0;
            operation_194_4372 <= 32'd0;
            operation_194_4384 <= 32'd0;
            operation_194_4386 <= 32'd0;
            operation_194_4388 <= 32'd0;
            operation_194_4390 <= 32'd0;
            operation_194_4392 <= 32'd0;
            operation_194_4394 <= 32'd0;
            operation_194_4396 <= 32'd0;
            operation_194_4398 <= 32'd0;
            operation_194_4400 <= 32'd0;
            operation_194_4402 <= 32'd0;
            operation_194_4414 <= 32'd0;
            operation_194_4416 <= 32'd0;
            operation_194_4418 <= 32'd0;
            operation_194_4420 <= 32'd0;
            operation_194_4422 <= 32'd0;
            operation_194_4424 <= 32'd0;
            operation_194_4426 <= 32'd0;
            operation_194_4428 <= 32'd0;
            operation_194_4430 <= 32'd0;
            operation_194_4432 <= 32'd0;
            operation_194_4444 <= 32'd0;
            operation_194_4445 <= 32'd0;
            operation_194_4447 <= 32'd0;
            operation_194_4448 <= 32'd0;
            operation_194_4450 <= 32'd0;
            operation_194_4451 <= 32'd0;
            operation_194_4453 <= 32'd0;
            operation_194_4454 <= 32'd0;
            operation_194_4456 <= 32'd0;
            operation_194_4457 <= 32'd0;
            operation_194_4459 <= 32'd0;
            operation_194_4460 <= 32'd0;
            operation_194_4462 <= 32'd0;
            operation_194_4463 <= 32'd0;
            operation_194_4465 <= 32'd0;
            operation_194_4466 <= 32'd0;
            operation_194_4468 <= 32'd0;
            operation_194_4470 <= 32'd0;
            operation_194_4473 <= 32'd0;
            operation_194_4474 <= 32'd0;
            operation_194_4475 <= 32'd0;
            operation_194_4477 <= 32'd0;
            operation_194_4478 <= 32'd0;
            operation_194_4479 <= 32'd0;
            operation_194_4481 <= 32'd0;
            operation_194_4482 <= 32'd0;
            operation_194_4483 <= 32'd0;
            operation_194_4485 <= 32'd0;
            operation_194_4486 <= 32'd0;
            operation_194_4487 <= 32'd0;
            operation_194_4489 <= 32'd0;
            operation_194_4490 <= 32'd0;
            operation_194_4491 <= 32'd0;
            operation_194_4493 <= 32'd0;
            operation_194_4494 <= 32'd0;
            operation_194_4495 <= 32'd0;
            operation_194_4497 <= 32'd0;
            operation_194_4498 <= 32'd0;
            operation_194_4499 <= 32'd0;
            operation_194_4501 <= 32'd0;
            operation_194_4502 <= 32'd0;
            operation_194_4503 <= 32'd0;
            operation_194_4506 <= 32'd0;
            operation_194_4507 <= 32'd0;
            operation_194_4509 <= 32'd0;
            operation_194_4510 <= 32'd0;
            operation_194_4512 <= 32'd0;
            operation_194_4513 <= 32'd0;
            operation_194_4515 <= 32'd0;
            operation_194_4516 <= 32'd0;
            operation_194_4518 <= 32'd0;
            operation_194_4519 <= 32'd0;
            operation_194_4521 <= 32'd0;
            operation_194_4522 <= 32'd0;
            operation_194_4524 <= 32'd0;
            operation_194_4525 <= 32'd0;
            operation_194_4527 <= 32'd0;
            operation_194_4528 <= 32'd0;
            operation_194_4530 <= 32'd0;
            operation_194_4532 <= 32'd0;
            operation_194_4537 <= 32'd0;
            operation_194_4538 <= 32'd0;
            operation_194_4539 <= 32'd0;
            operation_194_4541 <= 32'd0;
            operation_194_4542 <= 32'd0;
            operation_194_4543 <= 32'd0;
            operation_194_4545 <= 32'd0;
            operation_194_4546 <= 32'd0;
            operation_194_4547 <= 32'd0;
            operation_194_4549 <= 32'd0;
            operation_194_4550 <= 32'd0;
            operation_194_4551 <= 32'd0;
            operation_194_4553 <= 32'd0;
            operation_194_4554 <= 32'd0;
            operation_194_4555 <= 32'd0;
            operation_194_4557 <= 32'd0;
            operation_194_4558 <= 32'd0;
            operation_194_4559 <= 32'd0;
            operation_194_4561 <= 32'd0;
            operation_194_4562 <= 32'd0;
            operation_194_4563 <= 32'd0;
            operation_194_4565 <= 32'd0;
            operation_194_4566 <= 32'd0;
            operation_194_4567 <= 32'd0;
            operation_194_4571 <= 32'd0;
            operation_194_4574 <= 32'd0;
            operation_194_4577 <= 32'd0;
            operation_194_4580 <= 32'd0;
            operation_194_4582 <= 32'd0;
            operation_194_4584 <= 32'd0;
            operation_194_4586 <= 32'd0;
            operation_194_4588 <= 32'd0;
            operation_194_4590 <= 32'd0;
            operation_194_4596 <= 32'd0;
            operation_194_4597 <= 32'd0;
            operation_194_4598 <= 32'd0;
            operation_194_4599 <= 32'd0;
            operation_194_4601 <= 32'd0;
            operation_194_4603 <= 32'd0;
            operation_194_4605 <= 32'd0;
            operation_194_4607 <= 32'd0;
            operation_194_4609 <= 32'd0;
            operation_194_4611 <= 32'd0;
            operation_194_4613 <= 32'd0;
            operation_194_4615 <= 32'd0;
            operation_194_4617 <= 32'd0;
            operation_194_4619 <= 32'd0;
            operation_194_4621 <= 32'd0;
            operation_194_4631 <= 32'd0;
            operation_194_4632 <= 32'd0;
            operation_194_4633 <= 32'd0;
            operation_194_4634 <= 32'd0;
            operation_194_4646 <= 32'd0;
            operation_194_4648 <= 32'd0;
            operation_194_4663_latch <= 8'd0;
            operation_194_4664_latch <= 8'd0;
            operation_194_4673_latch <= 8'd0;
            operation_194_4674_latch <= 8'd0;
            operation_194_4675_latch <= 8'd0;
            operation_194_4676_latch <= 8'd0;
            operation_194_4677_latch <= 8'd0;
            operation_194_4678_latch <= 8'd0;
            operation_194_4679_latch <= 8'd0;
            operation_194_4680_latch <= 8'd0;
            operation_194_4681_latch <= 8'd0;
            operation_194_4682_latch <= 8'd0;
            operation_194_4683_latch <= 8'd0;
            operation_194_4684_latch <= 8'd0;
            operation_194_4685_latch <= 8'd0;
            operation_194_4686_latch <= 8'd0;
            operation_194_4687_latch <= 8'd0;
            operation_194_4688_latch <= 8'd0;
            operation_194_4689_latch <= 8'd0;
            operation_194_4690_latch <= 8'd0;
            operation_194_3845 <= 32'd0;
            operation_194_3849 <= 32'd0;
            operation_194_3851 <= 32'd0;
            operation_194_3853 <= 32'd0;
            operation_194_3855 <= 32'd0;
            operation_194_3857 <= 32'd0;
            operation_194_3859 <= 32'd0;
            operation_194_3861 <= 32'd0;
            operation_194_3863 <= 32'd0;
            operation_194_3875 <= 32'd0;
            operation_194_3877 <= 32'd0;
            operation_194_3879 <= 32'd0;
            operation_194_3881 <= 32'd0;
            operation_194_3883 <= 32'd0;
            operation_194_3885 <= 32'd0;
            operation_194_3887 <= 32'd0;
            operation_194_3889 <= 32'd0;
            operation_194_3891 <= 32'd0;
            operation_194_3893 <= 32'd0;
            operation_194_3895 <= 32'd0;
            operation_194_3897 <= 32'd0;
            operation_194_3899 <= 32'd0;
            operation_194_3901 <= 32'd0;
            operation_194_3903 <= 32'd0;
            operation_194_3905 <= 32'd0;
            operation_194_3925 <= 32'd0;
            operation_194_3927 <= 32'd0;
            operation_194_3929 <= 32'd0;
            operation_194_3931 <= 32'd0;
            operation_194_3933 <= 32'd0;
            operation_194_3935 <= 32'd0;
            operation_194_3937 <= 32'd0;
            operation_194_3939 <= 32'd0;
            operation_194_3941 <= 32'd0;
            operation_194_3943 <= 32'd0;
            operation_194_3955 <= 32'd0;
            operation_194_3957 <= 32'd0;
            operation_194_3959 <= 32'd0;
            operation_194_3961 <= 32'd0;
            operation_194_3963 <= 32'd0;
            operation_194_3965 <= 32'd0;
            operation_194_3967 <= 32'd0;
            operation_194_3969 <= 32'd0;
            operation_194_3971 <= 32'd0;
            operation_194_3973 <= 32'd0;
            operation_194_3985 <= 32'd0;
            operation_194_3987 <= 32'd0;
            operation_194_3989 <= 32'd0;
            operation_194_3991 <= 32'd0;
            operation_194_3993 <= 32'd0;
            operation_194_3995 <= 32'd0;
            operation_194_3997 <= 32'd0;
            operation_194_3999 <= 32'd0;
            operation_194_4001 <= 32'd0;
            operation_194_4003 <= 32'd0;
            operation_194_4015 <= 32'd0;
            operation_194_4016 <= 32'd0;
            operation_194_4018 <= 32'd0;
            operation_194_4019 <= 32'd0;
            operation_194_4021 <= 32'd0;
            operation_194_4022 <= 32'd0;
            operation_194_4024 <= 32'd0;
            operation_194_4025 <= 32'd0;
            operation_194_4027 <= 32'd0;
            operation_194_4028 <= 32'd0;
            operation_194_4030 <= 32'd0;
            operation_194_4031 <= 32'd0;
            operation_194_4033 <= 32'd0;
            operation_194_4034 <= 32'd0;
            operation_194_4036 <= 32'd0;
            operation_194_4037 <= 32'd0;
            operation_194_4039 <= 32'd0;
            operation_194_4041 <= 32'd0;
            operation_194_4044 <= 32'd0;
            operation_194_4045 <= 32'd0;
            operation_194_4046 <= 32'd0;
            operation_194_4048 <= 32'd0;
            operation_194_4049 <= 32'd0;
            operation_194_4050 <= 32'd0;
            operation_194_4052 <= 32'd0;
            operation_194_4053 <= 32'd0;
            operation_194_4054 <= 32'd0;
            operation_194_4056 <= 32'd0;
            operation_194_4057 <= 32'd0;
            operation_194_4058 <= 32'd0;
            operation_194_4060 <= 32'd0;
            operation_194_4061 <= 32'd0;
            operation_194_4062 <= 32'd0;
            operation_194_4064 <= 32'd0;
            operation_194_4065 <= 32'd0;
            operation_194_4066 <= 32'd0;
            operation_194_4068 <= 32'd0;
            operation_194_4069 <= 32'd0;
            operation_194_4070 <= 32'd0;
            operation_194_4072 <= 32'd0;
            operation_194_4073 <= 32'd0;
            operation_194_4074 <= 32'd0;
            operation_194_4077 <= 32'd0;
            operation_194_4078 <= 32'd0;
            operation_194_4080 <= 32'd0;
            operation_194_4081 <= 32'd0;
            operation_194_4083 <= 32'd0;
            operation_194_4084 <= 32'd0;
            operation_194_4086 <= 32'd0;
            operation_194_4087 <= 32'd0;
            operation_194_4089 <= 32'd0;
            operation_194_4090 <= 32'd0;
            operation_194_4092 <= 32'd0;
            operation_194_4093 <= 32'd0;
            operation_194_4095 <= 32'd0;
            operation_194_4096 <= 32'd0;
            operation_194_4098 <= 32'd0;
            operation_194_4099 <= 32'd0;
            operation_194_4101 <= 32'd0;
            operation_194_4103 <= 32'd0;
            operation_194_4108 <= 32'd0;
            operation_194_4109 <= 32'd0;
            operation_194_4110 <= 32'd0;
            operation_194_4112 <= 32'd0;
            operation_194_4113 <= 32'd0;
            operation_194_4114 <= 32'd0;
            operation_194_4116 <= 32'd0;
            operation_194_4117 <= 32'd0;
            operation_194_4118 <= 32'd0;
            operation_194_4120 <= 32'd0;
            operation_194_4121 <= 32'd0;
            operation_194_4122 <= 32'd0;
            operation_194_4124 <= 32'd0;
            operation_194_4125 <= 32'd0;
            operation_194_4126 <= 32'd0;
            operation_194_4128 <= 32'd0;
            operation_194_4129 <= 32'd0;
            operation_194_4130 <= 32'd0;
            operation_194_4132 <= 32'd0;
            operation_194_4133 <= 32'd0;
            operation_194_4134 <= 32'd0;
            operation_194_4136 <= 32'd0;
            operation_194_4137 <= 32'd0;
            operation_194_4138 <= 32'd0;
            operation_194_4142 <= 32'd0;
            operation_194_4145 <= 32'd0;
            operation_194_4148 <= 32'd0;
            operation_194_4151 <= 32'd0;
            operation_194_4153 <= 32'd0;
            operation_194_4155 <= 32'd0;
            operation_194_4157 <= 32'd0;
            operation_194_4159 <= 32'd0;
            operation_194_4161 <= 32'd0;
            operation_194_4167 <= 32'd0;
            operation_194_4168 <= 32'd0;
            operation_194_4169 <= 32'd0;
            operation_194_4170 <= 32'd0;
            operation_194_4172 <= 32'd0;
            operation_194_4174 <= 32'd0;
            operation_194_4176 <= 32'd0;
            operation_194_4178 <= 32'd0;
            operation_194_4180 <= 32'd0;
            operation_194_4182 <= 32'd0;
            operation_194_4184 <= 32'd0;
            operation_194_4186 <= 32'd0;
            operation_194_4188 <= 32'd0;
            operation_194_4190 <= 32'd0;
            operation_194_4192 <= 32'd0;
            operation_194_4202 <= 32'd0;
            operation_194_4203 <= 32'd0;
            operation_194_4204 <= 32'd0;
            operation_194_4205 <= 32'd0;
            operation_194_4217 <= 32'd0;
            operation_194_4219 <= 32'd0;
            operation_194_4234_latch <= 8'd0;
            operation_194_4235_latch <= 8'd0;
            operation_194_4244_latch <= 8'd0;
            operation_194_4245_latch <= 8'd0;
            operation_194_4246_latch <= 8'd0;
            operation_194_4247_latch <= 8'd0;
            operation_194_4248_latch <= 8'd0;
            operation_194_4249_latch <= 8'd0;
            operation_194_4250_latch <= 8'd0;
            operation_194_4251_latch <= 8'd0;
            operation_194_4252_latch <= 8'd0;
            operation_194_4253_latch <= 8'd0;
            operation_194_4254_latch <= 8'd0;
            operation_194_4255_latch <= 8'd0;
            operation_194_4256_latch <= 8'd0;
            operation_194_4257_latch <= 8'd0;
            operation_194_4258_latch <= 8'd0;
            operation_194_4259_latch <= 8'd0;
            operation_194_4260_latch <= 8'd0;
            operation_194_4261_latch <= 8'd0;
            operation_194_3416 <= 32'd0;
            operation_194_3420 <= 32'd0;
            operation_194_3422 <= 32'd0;
            operation_194_3424 <= 32'd0;
            operation_194_3426 <= 32'd0;
            operation_194_3428 <= 32'd0;
            operation_194_3430 <= 32'd0;
            operation_194_3432 <= 32'd0;
            operation_194_3434 <= 32'd0;
            operation_194_3446 <= 32'd0;
            operation_194_3448 <= 32'd0;
            operation_194_3450 <= 32'd0;
            operation_194_3452 <= 32'd0;
            operation_194_3454 <= 32'd0;
            operation_194_3456 <= 32'd0;
            operation_194_3458 <= 32'd0;
            operation_194_3460 <= 32'd0;
            operation_194_3462 <= 32'd0;
            operation_194_3464 <= 32'd0;
            operation_194_3466 <= 32'd0;
            operation_194_3468 <= 32'd0;
            operation_194_3470 <= 32'd0;
            operation_194_3472 <= 32'd0;
            operation_194_3474 <= 32'd0;
            operation_194_3476 <= 32'd0;
            operation_194_3496 <= 32'd0;
            operation_194_3498 <= 32'd0;
            operation_194_3500 <= 32'd0;
            operation_194_3502 <= 32'd0;
            operation_194_3504 <= 32'd0;
            operation_194_3506 <= 32'd0;
            operation_194_3508 <= 32'd0;
            operation_194_3510 <= 32'd0;
            operation_194_3512 <= 32'd0;
            operation_194_3514 <= 32'd0;
            operation_194_3526 <= 32'd0;
            operation_194_3528 <= 32'd0;
            operation_194_3530 <= 32'd0;
            operation_194_3532 <= 32'd0;
            operation_194_3534 <= 32'd0;
            operation_194_3536 <= 32'd0;
            operation_194_3538 <= 32'd0;
            operation_194_3540 <= 32'd0;
            operation_194_3542 <= 32'd0;
            operation_194_3544 <= 32'd0;
            operation_194_3556 <= 32'd0;
            operation_194_3558 <= 32'd0;
            operation_194_3560 <= 32'd0;
            operation_194_3562 <= 32'd0;
            operation_194_3564 <= 32'd0;
            operation_194_3566 <= 32'd0;
            operation_194_3568 <= 32'd0;
            operation_194_3570 <= 32'd0;
            operation_194_3572 <= 32'd0;
            operation_194_3574 <= 32'd0;
            operation_194_3586 <= 32'd0;
            operation_194_3587 <= 32'd0;
            operation_194_3589 <= 32'd0;
            operation_194_3590 <= 32'd0;
            operation_194_3592 <= 32'd0;
            operation_194_3593 <= 32'd0;
            operation_194_3595 <= 32'd0;
            operation_194_3596 <= 32'd0;
            operation_194_3598 <= 32'd0;
            operation_194_3599 <= 32'd0;
            operation_194_3601 <= 32'd0;
            operation_194_3602 <= 32'd0;
            operation_194_3604 <= 32'd0;
            operation_194_3605 <= 32'd0;
            operation_194_3607 <= 32'd0;
            operation_194_3608 <= 32'd0;
            operation_194_3610 <= 32'd0;
            operation_194_3612 <= 32'd0;
            operation_194_3615 <= 32'd0;
            operation_194_3616 <= 32'd0;
            operation_194_3617 <= 32'd0;
            operation_194_3619 <= 32'd0;
            operation_194_3620 <= 32'd0;
            operation_194_3621 <= 32'd0;
            operation_194_3623 <= 32'd0;
            operation_194_3624 <= 32'd0;
            operation_194_3625 <= 32'd0;
            operation_194_3627 <= 32'd0;
            operation_194_3628 <= 32'd0;
            operation_194_3629 <= 32'd0;
            operation_194_3631 <= 32'd0;
            operation_194_3632 <= 32'd0;
            operation_194_3633 <= 32'd0;
            operation_194_3635 <= 32'd0;
            operation_194_3636 <= 32'd0;
            operation_194_3637 <= 32'd0;
            operation_194_3639 <= 32'd0;
            operation_194_3640 <= 32'd0;
            operation_194_3641 <= 32'd0;
            operation_194_3643 <= 32'd0;
            operation_194_3644 <= 32'd0;
            operation_194_3645 <= 32'd0;
            operation_194_3648 <= 32'd0;
            operation_194_3649 <= 32'd0;
            operation_194_3651 <= 32'd0;
            operation_194_3652 <= 32'd0;
            operation_194_3654 <= 32'd0;
            operation_194_3655 <= 32'd0;
            operation_194_3657 <= 32'd0;
            operation_194_3658 <= 32'd0;
            operation_194_3660 <= 32'd0;
            operation_194_3661 <= 32'd0;
            operation_194_3663 <= 32'd0;
            operation_194_3664 <= 32'd0;
            operation_194_3666 <= 32'd0;
            operation_194_3667 <= 32'd0;
            operation_194_3669 <= 32'd0;
            operation_194_3670 <= 32'd0;
            operation_194_3672 <= 32'd0;
            operation_194_3674 <= 32'd0;
            operation_194_3679 <= 32'd0;
            operation_194_3680 <= 32'd0;
            operation_194_3681 <= 32'd0;
            operation_194_3683 <= 32'd0;
            operation_194_3684 <= 32'd0;
            operation_194_3685 <= 32'd0;
            operation_194_3687 <= 32'd0;
            operation_194_3688 <= 32'd0;
            operation_194_3689 <= 32'd0;
            operation_194_3691 <= 32'd0;
            operation_194_3692 <= 32'd0;
            operation_194_3693 <= 32'd0;
            operation_194_3695 <= 32'd0;
            operation_194_3696 <= 32'd0;
            operation_194_3697 <= 32'd0;
            operation_194_3699 <= 32'd0;
            operation_194_3700 <= 32'd0;
            operation_194_3701 <= 32'd0;
            operation_194_3703 <= 32'd0;
            operation_194_3704 <= 32'd0;
            operation_194_3705 <= 32'd0;
            operation_194_3707 <= 32'd0;
            operation_194_3708 <= 32'd0;
            operation_194_3709 <= 32'd0;
            operation_194_3713 <= 32'd0;
            operation_194_3716 <= 32'd0;
            operation_194_3719 <= 32'd0;
            operation_194_3722 <= 32'd0;
            operation_194_3724 <= 32'd0;
            operation_194_3726 <= 32'd0;
            operation_194_3728 <= 32'd0;
            operation_194_3730 <= 32'd0;
            operation_194_3732 <= 32'd0;
            operation_194_3738 <= 32'd0;
            operation_194_3739 <= 32'd0;
            operation_194_3740 <= 32'd0;
            operation_194_3741 <= 32'd0;
            operation_194_3743 <= 32'd0;
            operation_194_3745 <= 32'd0;
            operation_194_3747 <= 32'd0;
            operation_194_3749 <= 32'd0;
            operation_194_3751 <= 32'd0;
            operation_194_3753 <= 32'd0;
            operation_194_3755 <= 32'd0;
            operation_194_3757 <= 32'd0;
            operation_194_3759 <= 32'd0;
            operation_194_3761 <= 32'd0;
            operation_194_3763 <= 32'd0;
            operation_194_3773 <= 32'd0;
            operation_194_3774 <= 32'd0;
            operation_194_3775 <= 32'd0;
            operation_194_3776 <= 32'd0;
            operation_194_3788 <= 32'd0;
            operation_194_3790 <= 32'd0;
            operation_194_3805_latch <= 8'd0;
            operation_194_3806_latch <= 8'd0;
            operation_194_3815_latch <= 8'd0;
            operation_194_3816_latch <= 8'd0;
            operation_194_3817_latch <= 8'd0;
            operation_194_3818_latch <= 8'd0;
            operation_194_3819_latch <= 8'd0;
            operation_194_3820_latch <= 8'd0;
            operation_194_3821_latch <= 8'd0;
            operation_194_3822_latch <= 8'd0;
            operation_194_3823_latch <= 8'd0;
            operation_194_3824_latch <= 8'd0;
            operation_194_3825_latch <= 8'd0;
            operation_194_3826_latch <= 8'd0;
            operation_194_3827_latch <= 8'd0;
            operation_194_3828_latch <= 8'd0;
            operation_194_3829_latch <= 8'd0;
            operation_194_3830_latch <= 8'd0;
            operation_194_3831_latch <= 8'd0;
            operation_194_3832_latch <= 8'd0;
            operation_194_2987 <= 32'd0;
            operation_194_2991 <= 32'd0;
            operation_194_2993 <= 32'd0;
            operation_194_2995 <= 32'd0;
            operation_194_2997 <= 32'd0;
            operation_194_2999 <= 32'd0;
            operation_194_3001 <= 32'd0;
            operation_194_3003 <= 32'd0;
            operation_194_3005 <= 32'd0;
            operation_194_3017 <= 32'd0;
            operation_194_3019 <= 32'd0;
            operation_194_3021 <= 32'd0;
            operation_194_3023 <= 32'd0;
            operation_194_3025 <= 32'd0;
            operation_194_3027 <= 32'd0;
            operation_194_3029 <= 32'd0;
            operation_194_3031 <= 32'd0;
            operation_194_3033 <= 32'd0;
            operation_194_3035 <= 32'd0;
            operation_194_3037 <= 32'd0;
            operation_194_3039 <= 32'd0;
            operation_194_3041 <= 32'd0;
            operation_194_3043 <= 32'd0;
            operation_194_3045 <= 32'd0;
            operation_194_3047 <= 32'd0;
            operation_194_3067 <= 32'd0;
            operation_194_3069 <= 32'd0;
            operation_194_3071 <= 32'd0;
            operation_194_3073 <= 32'd0;
            operation_194_3075 <= 32'd0;
            operation_194_3077 <= 32'd0;
            operation_194_3079 <= 32'd0;
            operation_194_3081 <= 32'd0;
            operation_194_3083 <= 32'd0;
            operation_194_3085 <= 32'd0;
            operation_194_3097 <= 32'd0;
            operation_194_3099 <= 32'd0;
            operation_194_3101 <= 32'd0;
            operation_194_3103 <= 32'd0;
            operation_194_3105 <= 32'd0;
            operation_194_3107 <= 32'd0;
            operation_194_3109 <= 32'd0;
            operation_194_3111 <= 32'd0;
            operation_194_3113 <= 32'd0;
            operation_194_3115 <= 32'd0;
            operation_194_3127 <= 32'd0;
            operation_194_3129 <= 32'd0;
            operation_194_3131 <= 32'd0;
            operation_194_3133 <= 32'd0;
            operation_194_3135 <= 32'd0;
            operation_194_3137 <= 32'd0;
            operation_194_3139 <= 32'd0;
            operation_194_3141 <= 32'd0;
            operation_194_3143 <= 32'd0;
            operation_194_3145 <= 32'd0;
            operation_194_3157 <= 32'd0;
            operation_194_3158 <= 32'd0;
            operation_194_3160 <= 32'd0;
            operation_194_3161 <= 32'd0;
            operation_194_3163 <= 32'd0;
            operation_194_3164 <= 32'd0;
            operation_194_3166 <= 32'd0;
            operation_194_3167 <= 32'd0;
            operation_194_3169 <= 32'd0;
            operation_194_3170 <= 32'd0;
            operation_194_3172 <= 32'd0;
            operation_194_3173 <= 32'd0;
            operation_194_3175 <= 32'd0;
            operation_194_3176 <= 32'd0;
            operation_194_3178 <= 32'd0;
            operation_194_3179 <= 32'd0;
            operation_194_3181 <= 32'd0;
            operation_194_3183 <= 32'd0;
            operation_194_3186 <= 32'd0;
            operation_194_3187 <= 32'd0;
            operation_194_3188 <= 32'd0;
            operation_194_3190 <= 32'd0;
            operation_194_3191 <= 32'd0;
            operation_194_3192 <= 32'd0;
            operation_194_3194 <= 32'd0;
            operation_194_3195 <= 32'd0;
            operation_194_3196 <= 32'd0;
            operation_194_3198 <= 32'd0;
            operation_194_3199 <= 32'd0;
            operation_194_3200 <= 32'd0;
            operation_194_3202 <= 32'd0;
            operation_194_3203 <= 32'd0;
            operation_194_3204 <= 32'd0;
            operation_194_3206 <= 32'd0;
            operation_194_3207 <= 32'd0;
            operation_194_3208 <= 32'd0;
            operation_194_3210 <= 32'd0;
            operation_194_3211 <= 32'd0;
            operation_194_3212 <= 32'd0;
            operation_194_3214 <= 32'd0;
            operation_194_3215 <= 32'd0;
            operation_194_3216 <= 32'd0;
            operation_194_3219 <= 32'd0;
            operation_194_3220 <= 32'd0;
            operation_194_3222 <= 32'd0;
            operation_194_3223 <= 32'd0;
            operation_194_3225 <= 32'd0;
            operation_194_3226 <= 32'd0;
            operation_194_3228 <= 32'd0;
            operation_194_3229 <= 32'd0;
            operation_194_3231 <= 32'd0;
            operation_194_3232 <= 32'd0;
            operation_194_3234 <= 32'd0;
            operation_194_3235 <= 32'd0;
            operation_194_3237 <= 32'd0;
            operation_194_3238 <= 32'd0;
            operation_194_3240 <= 32'd0;
            operation_194_3241 <= 32'd0;
            operation_194_3243 <= 32'd0;
            operation_194_3245 <= 32'd0;
            operation_194_3250 <= 32'd0;
            operation_194_3251 <= 32'd0;
            operation_194_3252 <= 32'd0;
            operation_194_3254 <= 32'd0;
            operation_194_3255 <= 32'd0;
            operation_194_3256 <= 32'd0;
            operation_194_3258 <= 32'd0;
            operation_194_3259 <= 32'd0;
            operation_194_3260 <= 32'd0;
            operation_194_3262 <= 32'd0;
            operation_194_3263 <= 32'd0;
            operation_194_3264 <= 32'd0;
            operation_194_3266 <= 32'd0;
            operation_194_3267 <= 32'd0;
            operation_194_3268 <= 32'd0;
            operation_194_3270 <= 32'd0;
            operation_194_3271 <= 32'd0;
            operation_194_3272 <= 32'd0;
            operation_194_3274 <= 32'd0;
            operation_194_3275 <= 32'd0;
            operation_194_3276 <= 32'd0;
            operation_194_3278 <= 32'd0;
            operation_194_3279 <= 32'd0;
            operation_194_3280 <= 32'd0;
            operation_194_3284 <= 32'd0;
            operation_194_3287 <= 32'd0;
            operation_194_3290 <= 32'd0;
            operation_194_3293 <= 32'd0;
            operation_194_3295 <= 32'd0;
            operation_194_3297 <= 32'd0;
            operation_194_3299 <= 32'd0;
            operation_194_3301 <= 32'd0;
            operation_194_3303 <= 32'd0;
            operation_194_3309 <= 32'd0;
            operation_194_3310 <= 32'd0;
            operation_194_3311 <= 32'd0;
            operation_194_3312 <= 32'd0;
            operation_194_3314 <= 32'd0;
            operation_194_3316 <= 32'd0;
            operation_194_3318 <= 32'd0;
            operation_194_3320 <= 32'd0;
            operation_194_3322 <= 32'd0;
            operation_194_3324 <= 32'd0;
            operation_194_3326 <= 32'd0;
            operation_194_3328 <= 32'd0;
            operation_194_3330 <= 32'd0;
            operation_194_3332 <= 32'd0;
            operation_194_3334 <= 32'd0;
            operation_194_3344 <= 32'd0;
            operation_194_3345 <= 32'd0;
            operation_194_3346 <= 32'd0;
            operation_194_3347 <= 32'd0;
            operation_194_3359 <= 32'd0;
            operation_194_3361 <= 32'd0;
            operation_194_3376_latch <= 8'd0;
            operation_194_3377_latch <= 8'd0;
            operation_194_3386_latch <= 8'd0;
            operation_194_3387_latch <= 8'd0;
            operation_194_3388_latch <= 8'd0;
            operation_194_3389_latch <= 8'd0;
            operation_194_3390_latch <= 8'd0;
            operation_194_3391_latch <= 8'd0;
            operation_194_3392_latch <= 8'd0;
            operation_194_3393_latch <= 8'd0;
            operation_194_3394_latch <= 8'd0;
            operation_194_3395_latch <= 8'd0;
            operation_194_3396_latch <= 8'd0;
            operation_194_3397_latch <= 8'd0;
            operation_194_3398_latch <= 8'd0;
            operation_194_3399_latch <= 8'd0;
            operation_194_3400_latch <= 8'd0;
            operation_194_3401_latch <= 8'd0;
            operation_194_3402_latch <= 8'd0;
            operation_194_3403_latch <= 8'd0;
            operation_194_2558 <= 32'd0;
            operation_194_2562 <= 32'd0;
            operation_194_2564 <= 32'd0;
            operation_194_2566 <= 32'd0;
            operation_194_2568 <= 32'd0;
            operation_194_2570 <= 32'd0;
            operation_194_2572 <= 32'd0;
            operation_194_2574 <= 32'd0;
            operation_194_2576 <= 32'd0;
            operation_194_2588 <= 32'd0;
            operation_194_2590 <= 32'd0;
            operation_194_2592 <= 32'd0;
            operation_194_2594 <= 32'd0;
            operation_194_2596 <= 32'd0;
            operation_194_2598 <= 32'd0;
            operation_194_2600 <= 32'd0;
            operation_194_2602 <= 32'd0;
            operation_194_2604 <= 32'd0;
            operation_194_2606 <= 32'd0;
            operation_194_2608 <= 32'd0;
            operation_194_2610 <= 32'd0;
            operation_194_2612 <= 32'd0;
            operation_194_2614 <= 32'd0;
            operation_194_2616 <= 32'd0;
            operation_194_2618 <= 32'd0;
            operation_194_2638 <= 32'd0;
            operation_194_2640 <= 32'd0;
            operation_194_2642 <= 32'd0;
            operation_194_2644 <= 32'd0;
            operation_194_2646 <= 32'd0;
            operation_194_2648 <= 32'd0;
            operation_194_2650 <= 32'd0;
            operation_194_2652 <= 32'd0;
            operation_194_2654 <= 32'd0;
            operation_194_2656 <= 32'd0;
            operation_194_2668 <= 32'd0;
            operation_194_2670 <= 32'd0;
            operation_194_2672 <= 32'd0;
            operation_194_2674 <= 32'd0;
            operation_194_2676 <= 32'd0;
            operation_194_2678 <= 32'd0;
            operation_194_2680 <= 32'd0;
            operation_194_2682 <= 32'd0;
            operation_194_2684 <= 32'd0;
            operation_194_2686 <= 32'd0;
            operation_194_2698 <= 32'd0;
            operation_194_2700 <= 32'd0;
            operation_194_2702 <= 32'd0;
            operation_194_2704 <= 32'd0;
            operation_194_2706 <= 32'd0;
            operation_194_2708 <= 32'd0;
            operation_194_2710 <= 32'd0;
            operation_194_2712 <= 32'd0;
            operation_194_2714 <= 32'd0;
            operation_194_2716 <= 32'd0;
            operation_194_2728 <= 32'd0;
            operation_194_2729 <= 32'd0;
            operation_194_2731 <= 32'd0;
            operation_194_2732 <= 32'd0;
            operation_194_2734 <= 32'd0;
            operation_194_2735 <= 32'd0;
            operation_194_2737 <= 32'd0;
            operation_194_2738 <= 32'd0;
            operation_194_2740 <= 32'd0;
            operation_194_2741 <= 32'd0;
            operation_194_2743 <= 32'd0;
            operation_194_2744 <= 32'd0;
            operation_194_2746 <= 32'd0;
            operation_194_2747 <= 32'd0;
            operation_194_2749 <= 32'd0;
            operation_194_2750 <= 32'd0;
            operation_194_2752 <= 32'd0;
            operation_194_2754 <= 32'd0;
            operation_194_2757 <= 32'd0;
            operation_194_2758 <= 32'd0;
            operation_194_2759 <= 32'd0;
            operation_194_2761 <= 32'd0;
            operation_194_2762 <= 32'd0;
            operation_194_2763 <= 32'd0;
            operation_194_2765 <= 32'd0;
            operation_194_2766 <= 32'd0;
            operation_194_2767 <= 32'd0;
            operation_194_2769 <= 32'd0;
            operation_194_2770 <= 32'd0;
            operation_194_2771 <= 32'd0;
            operation_194_2773 <= 32'd0;
            operation_194_2774 <= 32'd0;
            operation_194_2775 <= 32'd0;
            operation_194_2777 <= 32'd0;
            operation_194_2778 <= 32'd0;
            operation_194_2779 <= 32'd0;
            operation_194_2781 <= 32'd0;
            operation_194_2782 <= 32'd0;
            operation_194_2783 <= 32'd0;
            operation_194_2785 <= 32'd0;
            operation_194_2786 <= 32'd0;
            operation_194_2787 <= 32'd0;
            operation_194_2790 <= 32'd0;
            operation_194_2791 <= 32'd0;
            operation_194_2793 <= 32'd0;
            operation_194_2794 <= 32'd0;
            operation_194_2796 <= 32'd0;
            operation_194_2797 <= 32'd0;
            operation_194_2799 <= 32'd0;
            operation_194_2800 <= 32'd0;
            operation_194_2802 <= 32'd0;
            operation_194_2803 <= 32'd0;
            operation_194_2805 <= 32'd0;
            operation_194_2806 <= 32'd0;
            operation_194_2808 <= 32'd0;
            operation_194_2809 <= 32'd0;
            operation_194_2811 <= 32'd0;
            operation_194_2812 <= 32'd0;
            operation_194_2814 <= 32'd0;
            operation_194_2816 <= 32'd0;
            operation_194_2821 <= 32'd0;
            operation_194_2822 <= 32'd0;
            operation_194_2823 <= 32'd0;
            operation_194_2825 <= 32'd0;
            operation_194_2826 <= 32'd0;
            operation_194_2827 <= 32'd0;
            operation_194_2829 <= 32'd0;
            operation_194_2830 <= 32'd0;
            operation_194_2831 <= 32'd0;
            operation_194_2833 <= 32'd0;
            operation_194_2834 <= 32'd0;
            operation_194_2835 <= 32'd0;
            operation_194_2837 <= 32'd0;
            operation_194_2838 <= 32'd0;
            operation_194_2839 <= 32'd0;
            operation_194_2841 <= 32'd0;
            operation_194_2842 <= 32'd0;
            operation_194_2843 <= 32'd0;
            operation_194_2845 <= 32'd0;
            operation_194_2846 <= 32'd0;
            operation_194_2847 <= 32'd0;
            operation_194_2849 <= 32'd0;
            operation_194_2850 <= 32'd0;
            operation_194_2851 <= 32'd0;
            operation_194_2855 <= 32'd0;
            operation_194_2858 <= 32'd0;
            operation_194_2861 <= 32'd0;
            operation_194_2864 <= 32'd0;
            operation_194_2866 <= 32'd0;
            operation_194_2868 <= 32'd0;
            operation_194_2870 <= 32'd0;
            operation_194_2872 <= 32'd0;
            operation_194_2874 <= 32'd0;
            operation_194_2880 <= 32'd0;
            operation_194_2881 <= 32'd0;
            operation_194_2882 <= 32'd0;
            operation_194_2883 <= 32'd0;
            operation_194_2885 <= 32'd0;
            operation_194_2887 <= 32'd0;
            operation_194_2889 <= 32'd0;
            operation_194_2891 <= 32'd0;
            operation_194_2893 <= 32'd0;
            operation_194_2895 <= 32'd0;
            operation_194_2897 <= 32'd0;
            operation_194_2899 <= 32'd0;
            operation_194_2901 <= 32'd0;
            operation_194_2903 <= 32'd0;
            operation_194_2905 <= 32'd0;
            operation_194_2915 <= 32'd0;
            operation_194_2916 <= 32'd0;
            operation_194_2917 <= 32'd0;
            operation_194_2918 <= 32'd0;
            operation_194_2930 <= 32'd0;
            operation_194_2932 <= 32'd0;
            operation_194_2947_latch <= 8'd0;
            operation_194_2948_latch <= 8'd0;
            operation_194_2957_latch <= 8'd0;
            operation_194_2958_latch <= 8'd0;
            operation_194_2959_latch <= 8'd0;
            operation_194_2960_latch <= 8'd0;
            operation_194_2961_latch <= 8'd0;
            operation_194_2962_latch <= 8'd0;
            operation_194_2963_latch <= 8'd0;
            operation_194_2964_latch <= 8'd0;
            operation_194_2965_latch <= 8'd0;
            operation_194_2966_latch <= 8'd0;
            operation_194_2967_latch <= 8'd0;
            operation_194_2968_latch <= 8'd0;
            operation_194_2969_latch <= 8'd0;
            operation_194_2970_latch <= 8'd0;
            operation_194_2971_latch <= 8'd0;
            operation_194_2972_latch <= 8'd0;
            operation_194_2973_latch <= 8'd0;
            operation_194_2974_latch <= 8'd0;
            operation_194_2129 <= 32'd0;
            operation_194_2133 <= 32'd0;
            operation_194_2135 <= 32'd0;
            operation_194_2137 <= 32'd0;
            operation_194_2139 <= 32'd0;
            operation_194_2141 <= 32'd0;
            operation_194_2143 <= 32'd0;
            operation_194_2145 <= 32'd0;
            operation_194_2147 <= 32'd0;
            operation_194_2159 <= 32'd0;
            operation_194_2161 <= 32'd0;
            operation_194_2163 <= 32'd0;
            operation_194_2165 <= 32'd0;
            operation_194_2167 <= 32'd0;
            operation_194_2169 <= 32'd0;
            operation_194_2171 <= 32'd0;
            operation_194_2173 <= 32'd0;
            operation_194_2175 <= 32'd0;
            operation_194_2177 <= 32'd0;
            operation_194_2179 <= 32'd0;
            operation_194_2181 <= 32'd0;
            operation_194_2183 <= 32'd0;
            operation_194_2185 <= 32'd0;
            operation_194_2187 <= 32'd0;
            operation_194_2189 <= 32'd0;
            operation_194_2209 <= 32'd0;
            operation_194_2211 <= 32'd0;
            operation_194_2213 <= 32'd0;
            operation_194_2215 <= 32'd0;
            operation_194_2217 <= 32'd0;
            operation_194_2219 <= 32'd0;
            operation_194_2221 <= 32'd0;
            operation_194_2223 <= 32'd0;
            operation_194_2225 <= 32'd0;
            operation_194_2227 <= 32'd0;
            operation_194_2239 <= 32'd0;
            operation_194_2241 <= 32'd0;
            operation_194_2243 <= 32'd0;
            operation_194_2245 <= 32'd0;
            operation_194_2247 <= 32'd0;
            operation_194_2249 <= 32'd0;
            operation_194_2251 <= 32'd0;
            operation_194_2253 <= 32'd0;
            operation_194_2255 <= 32'd0;
            operation_194_2257 <= 32'd0;
            operation_194_2269 <= 32'd0;
            operation_194_2271 <= 32'd0;
            operation_194_2273 <= 32'd0;
            operation_194_2275 <= 32'd0;
            operation_194_2277 <= 32'd0;
            operation_194_2279 <= 32'd0;
            operation_194_2281 <= 32'd0;
            operation_194_2283 <= 32'd0;
            operation_194_2285 <= 32'd0;
            operation_194_2287 <= 32'd0;
            operation_194_2299 <= 32'd0;
            operation_194_2300 <= 32'd0;
            operation_194_2302 <= 32'd0;
            operation_194_2303 <= 32'd0;
            operation_194_2305 <= 32'd0;
            operation_194_2306 <= 32'd0;
            operation_194_2308 <= 32'd0;
            operation_194_2309 <= 32'd0;
            operation_194_2311 <= 32'd0;
            operation_194_2312 <= 32'd0;
            operation_194_2314 <= 32'd0;
            operation_194_2315 <= 32'd0;
            operation_194_2317 <= 32'd0;
            operation_194_2318 <= 32'd0;
            operation_194_2320 <= 32'd0;
            operation_194_2321 <= 32'd0;
            operation_194_2323 <= 32'd0;
            operation_194_2325 <= 32'd0;
            operation_194_2328 <= 32'd0;
            operation_194_2329 <= 32'd0;
            operation_194_2330 <= 32'd0;
            operation_194_2332 <= 32'd0;
            operation_194_2333 <= 32'd0;
            operation_194_2334 <= 32'd0;
            operation_194_2336 <= 32'd0;
            operation_194_2337 <= 32'd0;
            operation_194_2338 <= 32'd0;
            operation_194_2340 <= 32'd0;
            operation_194_2341 <= 32'd0;
            operation_194_2342 <= 32'd0;
            operation_194_2344 <= 32'd0;
            operation_194_2345 <= 32'd0;
            operation_194_2346 <= 32'd0;
            operation_194_2348 <= 32'd0;
            operation_194_2349 <= 32'd0;
            operation_194_2350 <= 32'd0;
            operation_194_2352 <= 32'd0;
            operation_194_2353 <= 32'd0;
            operation_194_2354 <= 32'd0;
            operation_194_2356 <= 32'd0;
            operation_194_2357 <= 32'd0;
            operation_194_2358 <= 32'd0;
            operation_194_2361 <= 32'd0;
            operation_194_2362 <= 32'd0;
            operation_194_2364 <= 32'd0;
            operation_194_2365 <= 32'd0;
            operation_194_2367 <= 32'd0;
            operation_194_2368 <= 32'd0;
            operation_194_2370 <= 32'd0;
            operation_194_2371 <= 32'd0;
            operation_194_2373 <= 32'd0;
            operation_194_2374 <= 32'd0;
            operation_194_2376 <= 32'd0;
            operation_194_2377 <= 32'd0;
            operation_194_2379 <= 32'd0;
            operation_194_2380 <= 32'd0;
            operation_194_2382 <= 32'd0;
            operation_194_2383 <= 32'd0;
            operation_194_2385 <= 32'd0;
            operation_194_2387 <= 32'd0;
            operation_194_2392 <= 32'd0;
            operation_194_2393 <= 32'd0;
            operation_194_2394 <= 32'd0;
            operation_194_2396 <= 32'd0;
            operation_194_2397 <= 32'd0;
            operation_194_2398 <= 32'd0;
            operation_194_2400 <= 32'd0;
            operation_194_2401 <= 32'd0;
            operation_194_2402 <= 32'd0;
            operation_194_2404 <= 32'd0;
            operation_194_2405 <= 32'd0;
            operation_194_2406 <= 32'd0;
            operation_194_2408 <= 32'd0;
            operation_194_2409 <= 32'd0;
            operation_194_2410 <= 32'd0;
            operation_194_2412 <= 32'd0;
            operation_194_2413 <= 32'd0;
            operation_194_2414 <= 32'd0;
            operation_194_2416 <= 32'd0;
            operation_194_2417 <= 32'd0;
            operation_194_2418 <= 32'd0;
            operation_194_2420 <= 32'd0;
            operation_194_2421 <= 32'd0;
            operation_194_2422 <= 32'd0;
            operation_194_2426 <= 32'd0;
            operation_194_2429 <= 32'd0;
            operation_194_2432 <= 32'd0;
            operation_194_2435 <= 32'd0;
            operation_194_2437 <= 32'd0;
            operation_194_2439 <= 32'd0;
            operation_194_2441 <= 32'd0;
            operation_194_2443 <= 32'd0;
            operation_194_2445 <= 32'd0;
            operation_194_2451 <= 32'd0;
            operation_194_2452 <= 32'd0;
            operation_194_2453 <= 32'd0;
            operation_194_2454 <= 32'd0;
            operation_194_2456 <= 32'd0;
            operation_194_2458 <= 32'd0;
            operation_194_2460 <= 32'd0;
            operation_194_2462 <= 32'd0;
            operation_194_2464 <= 32'd0;
            operation_194_2466 <= 32'd0;
            operation_194_2468 <= 32'd0;
            operation_194_2470 <= 32'd0;
            operation_194_2472 <= 32'd0;
            operation_194_2474 <= 32'd0;
            operation_194_2476 <= 32'd0;
            operation_194_2486 <= 32'd0;
            operation_194_2487 <= 32'd0;
            operation_194_2488 <= 32'd0;
            operation_194_2489 <= 32'd0;
            operation_194_2501 <= 32'd0;
            operation_194_2503 <= 32'd0;
            operation_194_2518_latch <= 8'd0;
            operation_194_2519_latch <= 8'd0;
            operation_194_2528_latch <= 8'd0;
            operation_194_2529_latch <= 8'd0;
            operation_194_2530_latch <= 8'd0;
            operation_194_2531_latch <= 8'd0;
            operation_194_2532_latch <= 8'd0;
            operation_194_2533_latch <= 8'd0;
            operation_194_2534_latch <= 8'd0;
            operation_194_2535_latch <= 8'd0;
            operation_194_2536_latch <= 8'd0;
            operation_194_2537_latch <= 8'd0;
            operation_194_2538_latch <= 8'd0;
            operation_194_2539_latch <= 8'd0;
            operation_194_2540_latch <= 8'd0;
            operation_194_2541_latch <= 8'd0;
            operation_194_2542_latch <= 8'd0;
            operation_194_2543_latch <= 8'd0;
            operation_194_2544_latch <= 8'd0;
            operation_194_2545_latch <= 8'd0;
            operation_194_1700 <= 32'd0;
            operation_194_1704 <= 32'd0;
            operation_194_1706 <= 32'd0;
            operation_194_1708 <= 32'd0;
            operation_194_1710 <= 32'd0;
            operation_194_1712 <= 32'd0;
            operation_194_1714 <= 32'd0;
            operation_194_1716 <= 32'd0;
            operation_194_1718 <= 32'd0;
            operation_194_1730 <= 32'd0;
            operation_194_1732 <= 32'd0;
            operation_194_1734 <= 32'd0;
            operation_194_1736 <= 32'd0;
            operation_194_1738 <= 32'd0;
            operation_194_1740 <= 32'd0;
            operation_194_1742 <= 32'd0;
            operation_194_1744 <= 32'd0;
            operation_194_1746 <= 32'd0;
            operation_194_1748 <= 32'd0;
            operation_194_1750 <= 32'd0;
            operation_194_1752 <= 32'd0;
            operation_194_1754 <= 32'd0;
            operation_194_1756 <= 32'd0;
            operation_194_1758 <= 32'd0;
            operation_194_1760 <= 32'd0;
            operation_194_1780 <= 32'd0;
            operation_194_1782 <= 32'd0;
            operation_194_1784 <= 32'd0;
            operation_194_1786 <= 32'd0;
            operation_194_1788 <= 32'd0;
            operation_194_1790 <= 32'd0;
            operation_194_1792 <= 32'd0;
            operation_194_1794 <= 32'd0;
            operation_194_1796 <= 32'd0;
            operation_194_1798 <= 32'd0;
            operation_194_1810 <= 32'd0;
            operation_194_1812 <= 32'd0;
            operation_194_1814 <= 32'd0;
            operation_194_1816 <= 32'd0;
            operation_194_1818 <= 32'd0;
            operation_194_1820 <= 32'd0;
            operation_194_1822 <= 32'd0;
            operation_194_1824 <= 32'd0;
            operation_194_1826 <= 32'd0;
            operation_194_1828 <= 32'd0;
            operation_194_1840 <= 32'd0;
            operation_194_1842 <= 32'd0;
            operation_194_1844 <= 32'd0;
            operation_194_1846 <= 32'd0;
            operation_194_1848 <= 32'd0;
            operation_194_1850 <= 32'd0;
            operation_194_1852 <= 32'd0;
            operation_194_1854 <= 32'd0;
            operation_194_1856 <= 32'd0;
            operation_194_1858 <= 32'd0;
            operation_194_1870 <= 32'd0;
            operation_194_1871 <= 32'd0;
            operation_194_1873 <= 32'd0;
            operation_194_1874 <= 32'd0;
            operation_194_1876 <= 32'd0;
            operation_194_1877 <= 32'd0;
            operation_194_1879 <= 32'd0;
            operation_194_1880 <= 32'd0;
            operation_194_1882 <= 32'd0;
            operation_194_1883 <= 32'd0;
            operation_194_1885 <= 32'd0;
            operation_194_1886 <= 32'd0;
            operation_194_1888 <= 32'd0;
            operation_194_1889 <= 32'd0;
            operation_194_1891 <= 32'd0;
            operation_194_1892 <= 32'd0;
            operation_194_1894 <= 32'd0;
            operation_194_1896 <= 32'd0;
            operation_194_1899 <= 32'd0;
            operation_194_1900 <= 32'd0;
            operation_194_1901 <= 32'd0;
            operation_194_1903 <= 32'd0;
            operation_194_1904 <= 32'd0;
            operation_194_1905 <= 32'd0;
            operation_194_1907 <= 32'd0;
            operation_194_1908 <= 32'd0;
            operation_194_1909 <= 32'd0;
            operation_194_1911 <= 32'd0;
            operation_194_1912 <= 32'd0;
            operation_194_1913 <= 32'd0;
            operation_194_1915 <= 32'd0;
            operation_194_1916 <= 32'd0;
            operation_194_1917 <= 32'd0;
            operation_194_1919 <= 32'd0;
            operation_194_1920 <= 32'd0;
            operation_194_1921 <= 32'd0;
            operation_194_1923 <= 32'd0;
            operation_194_1924 <= 32'd0;
            operation_194_1925 <= 32'd0;
            operation_194_1927 <= 32'd0;
            operation_194_1928 <= 32'd0;
            operation_194_1929 <= 32'd0;
            operation_194_1932 <= 32'd0;
            operation_194_1933 <= 32'd0;
            operation_194_1935 <= 32'd0;
            operation_194_1936 <= 32'd0;
            operation_194_1938 <= 32'd0;
            operation_194_1939 <= 32'd0;
            operation_194_1941 <= 32'd0;
            operation_194_1942 <= 32'd0;
            operation_194_1944 <= 32'd0;
            operation_194_1945 <= 32'd0;
            operation_194_1947 <= 32'd0;
            operation_194_1948 <= 32'd0;
            operation_194_1950 <= 32'd0;
            operation_194_1951 <= 32'd0;
            operation_194_1953 <= 32'd0;
            operation_194_1954 <= 32'd0;
            operation_194_1956 <= 32'd0;
            operation_194_1958 <= 32'd0;
            operation_194_1963 <= 32'd0;
            operation_194_1964 <= 32'd0;
            operation_194_1965 <= 32'd0;
            operation_194_1967 <= 32'd0;
            operation_194_1968 <= 32'd0;
            operation_194_1969 <= 32'd0;
            operation_194_1971 <= 32'd0;
            operation_194_1972 <= 32'd0;
            operation_194_1973 <= 32'd0;
            operation_194_1975 <= 32'd0;
            operation_194_1976 <= 32'd0;
            operation_194_1977 <= 32'd0;
            operation_194_1979 <= 32'd0;
            operation_194_1980 <= 32'd0;
            operation_194_1981 <= 32'd0;
            operation_194_1983 <= 32'd0;
            operation_194_1984 <= 32'd0;
            operation_194_1985 <= 32'd0;
            operation_194_1987 <= 32'd0;
            operation_194_1988 <= 32'd0;
            operation_194_1989 <= 32'd0;
            operation_194_1991 <= 32'd0;
            operation_194_1992 <= 32'd0;
            operation_194_1993 <= 32'd0;
            operation_194_1997 <= 32'd0;
            operation_194_2000 <= 32'd0;
            operation_194_2003 <= 32'd0;
            operation_194_2006 <= 32'd0;
            operation_194_2008 <= 32'd0;
            operation_194_2010 <= 32'd0;
            operation_194_2012 <= 32'd0;
            operation_194_2014 <= 32'd0;
            operation_194_2016 <= 32'd0;
            operation_194_2022 <= 32'd0;
            operation_194_2023 <= 32'd0;
            operation_194_2024 <= 32'd0;
            operation_194_2025 <= 32'd0;
            operation_194_2027 <= 32'd0;
            operation_194_2029 <= 32'd0;
            operation_194_2031 <= 32'd0;
            operation_194_2033 <= 32'd0;
            operation_194_2035 <= 32'd0;
            operation_194_2037 <= 32'd0;
            operation_194_2039 <= 32'd0;
            operation_194_2041 <= 32'd0;
            operation_194_2043 <= 32'd0;
            operation_194_2045 <= 32'd0;
            operation_194_2047 <= 32'd0;
            operation_194_2057 <= 32'd0;
            operation_194_2058 <= 32'd0;
            operation_194_2059 <= 32'd0;
            operation_194_2060 <= 32'd0;
            operation_194_2072 <= 32'd0;
            operation_194_2074 <= 32'd0;
            operation_194_2089_latch <= 8'd0;
            operation_194_2090_latch <= 8'd0;
            operation_194_2099_latch <= 8'd0;
            operation_194_2100_latch <= 8'd0;
            operation_194_2101_latch <= 8'd0;
            operation_194_2102_latch <= 8'd0;
            operation_194_2103_latch <= 8'd0;
            operation_194_2104_latch <= 8'd0;
            operation_194_2105_latch <= 8'd0;
            operation_194_2106_latch <= 8'd0;
            operation_194_2107_latch <= 8'd0;
            operation_194_2108_latch <= 8'd0;
            operation_194_2109_latch <= 8'd0;
            operation_194_2110_latch <= 8'd0;
            operation_194_2111_latch <= 8'd0;
            operation_194_2112_latch <= 8'd0;
            operation_194_2113_latch <= 8'd0;
            operation_194_2114_latch <= 8'd0;
            operation_194_2115_latch <= 8'd0;
            operation_194_2116_latch <= 8'd0;
            operation_194_126 <= 32'd0;
            operation_194_6 <= 32'd0;
            operation_194_22 <= 32'd0;
            operation_194_38 <= 32'd0;
            operation_194_54 <= 32'd0;
            operation_194_70 <= 32'd0;
            operation_194_86 <= 32'd0;
            operation_194_102 <= 32'd0;
            operation_194_118 <= 32'd0;
            operation_194_14 <= 32'd0;
            operation_194_30 <= 32'd0;
            operation_194_46 <= 32'd0;
            operation_194_62 <= 32'd0;
            operation_194_78 <= 32'd0;
            operation_194_94 <= 32'd0;
            operation_194_110 <= 32'd0;
            control_194_follow <= 1'd0;
            control_194_start <= 1'd0;
            control_194_83 <= 1'd0;
            control_194_82 <= 1'd0;
            control_194_81 <= 1'd0;
            control_194_80 <= 1'd0;
            control_194_79 <= 1'd0;
            control_194_78 <= 1'd0;
            control_194_77 <= 1'd0;
            control_194_76 <= 1'd0;
            control_194_75 <= 1'd0;
            control_194_74 <= 1'd0;
            control_194_73 <= 1'd0;
            control_194_72 <= 1'd0;
            control_194_71 <= 1'd0;
            control_194_70 <= 1'd0;
            control_194_69 <= 1'd0;
            control_194_68 <= 1'd0;
            control_194_67 <= 1'd0;
            control_194_66 <= 1'd0;
            control_194_65 <= 1'd0;
            control_194_64 <= 1'd0;
            control_194_63 <= 1'd0;
            control_194_62 <= 1'd0;
            control_194_61 <= 1'd0;
            control_194_60 <= 1'd0;
            control_194_59 <= 1'd0;
            control_194_58 <= 1'd0;
            control_194_57 <= 1'd0;
            control_194_56 <= 1'd0;
            control_194_55 <= 1'd0;
            control_194_54 <= 1'd0;
            control_194_53 <= 1'd0;
            control_194_52 <= 1'd0;
            control_194_51 <= 1'd0;
            control_194_50 <= 1'd0;
            control_194_49 <= 1'd0;
            control_194_48 <= 1'd0;
            control_194_47 <= 1'd0;
            control_194_46 <= 1'd0;
            control_194_45 <= 1'd0;
            control_194_44 <= 1'd0;
            control_194_43 <= 1'd0;
            control_194_42 <= 1'd0;
            control_194_41 <= 1'd0;
            control_194_40 <= 1'd0;
            control_194_39 <= 1'd0;
            control_194_38 <= 1'd0;
            control_194_37 <= 1'd0;
            control_194_36 <= 1'd0;
            control_194_35 <= 1'd0;
            control_194_34 <= 1'd0;
            control_194_33 <= 1'd0;
            control_194_32 <= 1'd0;
            control_194_31 <= 1'd0;
            control_194_30 <= 1'd0;
            control_194_29 <= 1'd0;
            control_194_28 <= 1'd0;
            control_194_27 <= 1'd0;
            control_194_26 <= 1'd0;
            control_194_25 <= 1'd0;
            control_194_24 <= 1'd0;
            control_194_23 <= 1'd0;
            control_194_22 <= 1'd0;
            control_194_21 <= 1'd0;
            control_194_20 <= 1'd0;
            control_194_19 <= 1'd0;
            control_194_18 <= 1'd0;
            control_194_17 <= 1'd0;
            control_194_16 <= 1'd0;
            control_194_15 <= 1'd0;
            control_194_14 <= 1'd0;
            control_194_13 <= 1'd0;
            control_194_12 <= 1'd0;
            control_194_11 <= 1'd0;
            control_194_10 <= 1'd0;
            control_194_9 <= 1'd0;
            control_194_8 <= 1'd0;
            control_194_7 <= 1'd0;
            control_194_6 <= 1'd0;
            control_194_5 <= 1'd0;
            control_194_4 <= 1'd0;
            control_194_3 <= 1'd0;
            control_194_2 <= 1'd0;
            control_194_1 <= 1'd0;
            input_key_194_follow <= 128'd0;
            input_in_194_follow <= 128'd0;
            lookup_sbox_0_output <= 8'd0;
            lookup_sbox_1_output <= 8'd0;
            lookup_sbox_2_output <= 8'd0;
            lookup_sbox_3_output <= 8'd0;
            lookup_sbox_4_output <= 8'd0;
            lookup_sbox_5_output <= 8'd0;
            lookup_sbox_6_output <= 8'd0;
            lookup_sbox_7_output <= 8'd0;
            lookup_sbox_8_output <= 8'd0;
            lookup_sbox_9_output <= 8'd0;
            lookup_sbox_10_output <= 8'd0;
            lookup_sbox_11_output <= 8'd0;
            lookup_sbox_12_output <= 8'd0;
            lookup_sbox_13_output <= 8'd0;
            lookup_sbox_14_output <= 8'd0;
            lookup_sbox_15_output <= 8'd0;
            lookup_sbox_16_output <= 8'd0;
            lookup_sbox_17_output <= 8'd0;
            lookup_sbox_18_output <= 8'd0;
            lookup_sbox_19_output <= 8'd0;
            lookup_sbox_20_output <= 8'd0;
            lookup_sbox_21_output <= 8'd0;
            lookup_sbox_22_output <= 8'd0;
            lookup_sbox_23_output <= 8'd0;
            lookup_sbox_24_output <= 8'd0;
            lookup_sbox_25_output <= 8'd0;
            lookup_sbox_26_output <= 8'd0;
            lookup_sbox_27_output <= 8'd0;
            lookup_sbox_28_output <= 8'd0;
            lookup_sbox_29_output <= 8'd0;
            lookup_sbox_30_output <= 8'd0;
            lookup_sbox_31_output <= 8'd0;
            startfollow <= 1'd0;
        end
    else
        begin
            AES128_encrypt <= ((control_194_follow)?(return_194):(AES128_encrypt));
            finish <= ((!((start)&&(!(startfollow))))&&((finish)||(control_194_end)));
            control_194_start <= ((start)&&(!(startfollow)));
            operation_194_1664 <= ((operation_194_1661)^(operation_194_1663));
            operation_194_1536 <= ((operation_194_5133)^(operation_194_1535));
            operation_194_1680 <= ((operation_194_1677)^(operation_194_1679));
            operation_194_1632 <= ((operation_194_1629)^(operation_194_1535));
            operation_194_1672 <= ((operation_194_1669)^(operation_194_1671));
            operation_194_1688 <= ((operation_194_1685)^(operation_194_1687));
            operation_194_1504 <= ((operation_194_5160)^(operation_194_1503));
            operation_194_1552 <= ((operation_194_5151)^(operation_194_1551));
            operation_194_1648 <= ((operation_194_1645)^(operation_194_1551));
            operation_194_1600 <= ((operation_194_1597)^(operation_194_1503));
            operation_194_1544 <= ((operation_194_5195)^(operation_194_1543));
            operation_194_1560 <= ((operation_194_5193)^(operation_194_1559));
            operation_194_1656 <= ((operation_194_1653)^(operation_194_1559));
            operation_194_1640 <= ((operation_194_1637)^(operation_194_1543));
            operation_194_1472 <= ((operation_194_5232)^(operation_194_1471));
            operation_194_1520 <= ((operation_194_5231)^(operation_194_1519));
            operation_194_1616 <= ((operation_194_1613)^(operation_194_1519));
            operation_194_1568 <= ((operation_194_1565)^(operation_194_1471));
            operation_194_1512 <= ((operation_194_5262)^(operation_194_1511));
            operation_194_1528 <= ((operation_194_5261)^(operation_194_1527));
            operation_194_1624 <= ((operation_194_1621)^(operation_194_1527));
            operation_194_1608 <= ((operation_194_1605)^(operation_194_1511));
            operation_194_1440 <= ((operation_194_5292)^(operation_194_1439));
            operation_194_1488 <= ((operation_194_5291)^(operation_194_1487));
            operation_194_1584 <= ((operation_194_1581)^(operation_194_1487));
            operation_194_1432 <= ((operation_194_1428)^(operation_194_5601));
            operation_194_1480 <= ((operation_194_5330)^(operation_194_1479));
            operation_194_1496 <= ((operation_194_5329)^(operation_194_1495));
            operation_194_1592 <= ((operation_194_1589)^(operation_194_1495));
            operation_194_1576 <= ((operation_194_1573)^(operation_194_1479));
            operation_194_1456 <= ((operation_194_5391)^(operation_194_1455));
            operation_194_1448 <= ((operation_194_5450)^(operation_194_1447));
            operation_194_1464 <= ((operation_194_5449)^(operation_194_1463));
            operation_194_1338_latch <= (operation_194_1338);
            operation_194_1328_latch <= (operation_194_1328);
            operation_194_1318_latch <= (operation_194_1318);
            operation_194_1308_latch <= (operation_194_1308);
            operation_194_1298_latch <= (operation_194_1298);
            operation_194_1288_latch <= (operation_194_1288);
            operation_194_1278_latch <= (operation_194_1278);
            operation_194_1268_latch <= (operation_194_1268);
            operation_194_1273_latch <= (operation_194_1273);
            operation_194_1283_latch <= (operation_194_1283);
            operation_194_1293_latch <= (operation_194_1293);
            operation_194_1303_latch <= (operation_194_1303);
            operation_194_1313_latch <= (operation_194_1313);
            operation_194_1323_latch <= (operation_194_1323);
            operation_194_1333_latch <= (operation_194_1333);
            operation_194_1343_latch <= (operation_194_1343);
            operation_194_1413_latch <= (operation_194_1413);
            operation_194_1423_latch <= (operation_194_1423);
            operation_194_1408_latch <= (operation_194_1408);
            operation_194_1418_latch <= (operation_194_1418);
            operation_194_5132 <= ((operation_194_5153)^(operation_194_5133));
            operation_194_5136 <= ((operation_194_4704)^(operation_194_5160));
            operation_194_5138 <= ((operation_194_5159)^(operation_194_5292));
            operation_194_5140 <= ((operation_194_5158)^(operation_194_5391));
            operation_194_5142 <= ((operation_194_5157)^(operation_194_5232));
            operation_194_5144 <= ((operation_194_5156)^(operation_194_5291));
            operation_194_5146 <= ((operation_194_5155)^(operation_194_5160));
            operation_194_5148 <= ((operation_194_5154)^(operation_194_5231));
            operation_194_5150 <= ((operation_194_5152)^(operation_194_5151));
            operation_194_5162 <= ((operation_194_5499)^(operation_194_5210));
            operation_194_5164 <= ((operation_194_5500)^(operation_194_5209));
            operation_194_5166 <= ((operation_194_5497)^(operation_194_5208));
            operation_194_5168 <= ((operation_194_5498)^(operation_194_5207));
            operation_194_5170 <= ((operation_194_5495)^(operation_194_5206));
            operation_194_5172 <= ((operation_194_5496)^(operation_194_5205));
            operation_194_5174 <= ((operation_194_5493)^(operation_194_5204));
            operation_194_5176 <= ((operation_194_5494)^(operation_194_5203));
            operation_194_5178 <= ((operation_194_5202)^(operation_194_5450));
            operation_194_5180 <= ((operation_194_5201)^(operation_194_5449));
            operation_194_5182 <= ((operation_194_5200)^(operation_194_5330));
            operation_194_5184 <= ((operation_194_5199)^(operation_194_5329));
            operation_194_5186 <= ((operation_194_5198)^(operation_194_5262));
            operation_194_5188 <= ((operation_194_5197)^(operation_194_5261));
            operation_194_5190 <= ((operation_194_5196)^(operation_194_5195));
            operation_194_5192 <= ((operation_194_5194)^(operation_194_5193));
            operation_194_5212 <= ((operation_194_5530)^(operation_194_5240));
            operation_194_5214 <= ((operation_194_5529)^(operation_194_5239));
            operation_194_5216 <= ((operation_194_5528)^(operation_194_5238));
            operation_194_5218 <= ((operation_194_5527)^(operation_194_5237));
            operation_194_5220 <= ((operation_194_5526)^(operation_194_5236));
            operation_194_5222 <= ((operation_194_5525)^(operation_194_5235));
            operation_194_5224 <= ((operation_194_5524)^(operation_194_5234));
            operation_194_5226 <= ((operation_194_5523)^(operation_194_5233));
            operation_194_5228 <= ((operation_194_4731)^(operation_194_5232));
            operation_194_5230 <= ((operation_194_4722)^(operation_194_5231));
            operation_194_5242 <= ((operation_194_5270)^(operation_194_5394));
            operation_194_5244 <= ((operation_194_5269)^(operation_194_5394));
            operation_194_5246 <= ((operation_194_5268)^(operation_194_5453));
            operation_194_5248 <= ((operation_194_5267)^(operation_194_5453));
            operation_194_5250 <= ((operation_194_5266)^(operation_194_5393));
            operation_194_5252 <= ((operation_194_5265)^(operation_194_5393));
            operation_194_5254 <= ((operation_194_5264)^(operation_194_5452));
            operation_194_5256 <= ((operation_194_5263)^(operation_194_5452));
            operation_194_5258 <= ((operation_194_4766)^(operation_194_5262));
            operation_194_5260 <= ((operation_194_4764)^(operation_194_5261));
            operation_194_5272 <= ((operation_194_5300)^(operation_194_5394));
            operation_194_5274 <= ((operation_194_5299)^(operation_194_5394));
            operation_194_5276 <= ((operation_194_5298)^(operation_194_5453));
            operation_194_5278 <= ((operation_194_5297)^(operation_194_5453));
            operation_194_5280 <= ((operation_194_5296)^(operation_194_5393));
            operation_194_5282 <= ((operation_194_5295)^(operation_194_5393));
            operation_194_5284 <= ((operation_194_5294)^(operation_194_5452));
            operation_194_5286 <= ((operation_194_5293)^(operation_194_5452));
            operation_194_5288 <= ((operation_194_4803)^(operation_194_5292));
            operation_194_5290 <= ((operation_194_4802)^(operation_194_5291));
            operation_194_5302 <= ((operation_194_5361)^(operation_194_5303));
            operation_194_5303 <= ((operation_194_5359)*(operation_194_5597));
            operation_194_5305 <= ((operation_194_5357)^(operation_194_5306));
            operation_194_5306 <= ((operation_194_5355)*(operation_194_5597));
            operation_194_5308 <= ((operation_194_5353)^(operation_194_5309));
            operation_194_5309 <= ((operation_194_5351)*(operation_194_5597));
            operation_194_5311 <= ((operation_194_5349)^(operation_194_5312));
            operation_194_5312 <= ((operation_194_5347)*(operation_194_5597));
            operation_194_5314 <= ((operation_194_5345)^(operation_194_5315));
            operation_194_5315 <= ((operation_194_5343)*(operation_194_5597));
            operation_194_5317 <= ((operation_194_5341)^(operation_194_5318));
            operation_194_5318 <= ((operation_194_5339)*(operation_194_5597));
            operation_194_5320 <= ((operation_194_5337)^(operation_194_5321));
            operation_194_5321 <= ((operation_194_5335)*(operation_194_5597));
            operation_194_5323 <= ((operation_194_5333)^(operation_194_5324));
            operation_194_5324 <= ((operation_194_5331)*(operation_194_5597));
            operation_194_5326 <= ((operation_194_4833)^(operation_194_5330));
            operation_194_5328 <= ((operation_194_4832)^(operation_194_5329));
            operation_194_5331 <= ((operation_194_5332)&(operation_194_5557));
            operation_194_5332 <= ((operation_194_5334)>>(operation_194_2119));
            operation_194_5333 <= ((operation_194_5334)<<(operation_194_5557));
            operation_194_5335 <= ((operation_194_5336)&(operation_194_5557));
            operation_194_5336 <= ((operation_194_5338)>>(operation_194_2119));
            operation_194_5337 <= ((operation_194_5338)<<(operation_194_5557));
            operation_194_5339 <= ((operation_194_5340)&(operation_194_5557));
            operation_194_5340 <= ((operation_194_5342)>>(operation_194_2119));
            operation_194_5341 <= ((operation_194_5342)<<(operation_194_5557));
            operation_194_5343 <= ((operation_194_5344)&(operation_194_5557));
            operation_194_5344 <= ((operation_194_5346)>>(operation_194_2119));
            operation_194_5345 <= ((operation_194_5346)<<(operation_194_5557));
            operation_194_5347 <= ((operation_194_5348)&(operation_194_5557));
            operation_194_5348 <= ((operation_194_5350)>>(operation_194_2119));
            operation_194_5349 <= ((operation_194_5350)<<(operation_194_5557));
            operation_194_5351 <= ((operation_194_5352)&(operation_194_5557));
            operation_194_5352 <= ((operation_194_5354)>>(operation_194_2119));
            operation_194_5353 <= ((operation_194_5354)<<(operation_194_5557));
            operation_194_5355 <= ((operation_194_5356)&(operation_194_5557));
            operation_194_5356 <= ((operation_194_5358)>>(operation_194_2119));
            operation_194_5357 <= ((operation_194_5358)<<(operation_194_5557));
            operation_194_5359 <= ((operation_194_5360)&(operation_194_5557));
            operation_194_5360 <= ((operation_194_5362)>>(operation_194_2119));
            operation_194_5361 <= ((operation_194_5362)<<(operation_194_5557));
            operation_194_5364 <= ((operation_194_5425)^(operation_194_5365));
            operation_194_5365 <= ((operation_194_5423)*(operation_194_5597));
            operation_194_5367 <= ((operation_194_5421)^(operation_194_5368));
            operation_194_5368 <= ((operation_194_5419)*(operation_194_5597));
            operation_194_5370 <= ((operation_194_5417)^(operation_194_5371));
            operation_194_5371 <= ((operation_194_5415)*(operation_194_5597));
            operation_194_5373 <= ((operation_194_5413)^(operation_194_5374));
            operation_194_5374 <= ((operation_194_5411)*(operation_194_5597));
            operation_194_5376 <= ((operation_194_5409)^(operation_194_5377));
            operation_194_5377 <= ((operation_194_5407)*(operation_194_5597));
            operation_194_5379 <= ((operation_194_5405)^(operation_194_5380));
            operation_194_5380 <= ((operation_194_5403)*(operation_194_5597));
            operation_194_5382 <= ((operation_194_5401)^(operation_194_5383));
            operation_194_5383 <= ((operation_194_5399)*(operation_194_5597));
            operation_194_5385 <= ((operation_194_5397)^(operation_194_5386));
            operation_194_5386 <= ((operation_194_5395)*(operation_194_5597));
            operation_194_5388 <= ((operation_194_4863)^(operation_194_5392));
            operation_194_5390 <= ((operation_194_4862)^(operation_194_5391));
            operation_194_5395 <= ((operation_194_5396)&(operation_194_5557));
            operation_194_5396 <= ((operation_194_5398)>>(operation_194_2119));
            operation_194_5397 <= ((operation_194_5398)<<(operation_194_5557));
            operation_194_5399 <= ((operation_194_5400)&(operation_194_5557));
            operation_194_5400 <= ((operation_194_5402)>>(operation_194_2119));
            operation_194_5401 <= ((operation_194_5402)<<(operation_194_5557));
            operation_194_5403 <= ((operation_194_5404)&(operation_194_5557));
            operation_194_5404 <= ((operation_194_5406)>>(operation_194_2119));
            operation_194_5405 <= ((operation_194_5406)<<(operation_194_5557));
            operation_194_5407 <= ((operation_194_5408)&(operation_194_5557));
            operation_194_5408 <= ((operation_194_5410)>>(operation_194_2119));
            operation_194_5409 <= ((operation_194_5410)<<(operation_194_5557));
            operation_194_5411 <= ((operation_194_5412)&(operation_194_5557));
            operation_194_5412 <= ((operation_194_5414)>>(operation_194_2119));
            operation_194_5413 <= ((operation_194_5414)<<(operation_194_5557));
            operation_194_5415 <= ((operation_194_5416)&(operation_194_5557));
            operation_194_5416 <= ((operation_194_5418)>>(operation_194_2119));
            operation_194_5417 <= ((operation_194_5418)<<(operation_194_5557));
            operation_194_5419 <= ((operation_194_5420)&(operation_194_5557));
            operation_194_5420 <= ((operation_194_5422)>>(operation_194_2119));
            operation_194_5421 <= ((operation_194_5422)<<(operation_194_5557));
            operation_194_5423 <= ((operation_194_5424)&(operation_194_5557));
            operation_194_5424 <= ((operation_194_5426)>>(operation_194_2119));
            operation_194_5425 <= ((operation_194_5426)<<(operation_194_5557));
            operation_194_5429 <= ((operation_194_5500)^(operation_194_5529));
            operation_194_5432 <= ((operation_194_5498)^(operation_194_5527));
            operation_194_5435 <= ((operation_194_5496)^(operation_194_5525));
            operation_194_5438 <= ((operation_194_5494)^(operation_194_5523));
            operation_194_5440 <= ((operation_194_5456)^(operation_194_5529));
            operation_194_5442 <= ((operation_194_5454)^(operation_194_5525));
            operation_194_5444 <= ((operation_194_5451)^(operation_194_5597));
            operation_194_5446 <= ((operation_194_4901)^(operation_194_5450));
            operation_194_5448 <= ((operation_194_4900)^(operation_194_5449));
            operation_194_5454 <= ((operation_194_5455)^(operation_194_5496));
            operation_194_5455 <= ((operation_194_5495)^(operation_194_5526));
            operation_194_5456 <= ((operation_194_5457)^(operation_194_5500));
            operation_194_5457 <= ((operation_194_5499)^(operation_194_5530));
            operation_194_5459 <= ((operation_194_5530)^(operation_194_5500));
            operation_194_5461 <= ((operation_194_5529)^(operation_194_5499));
            operation_194_5463 <= ((operation_194_5528)^(operation_194_5498));
            operation_194_5465 <= ((operation_194_5527)^(operation_194_5497));
            operation_194_5467 <= ((operation_194_5526)^(operation_194_5496));
            operation_194_5469 <= ((operation_194_5525)^(operation_194_5495));
            operation_194_5471 <= ((operation_194_5524)^(operation_194_5494));
            operation_194_5473 <= ((operation_194_5523)^(operation_194_5493));
            operation_194_5475 <= ((operation_194_5491)^(operation_194_5527));
            operation_194_5477 <= ((operation_194_5489)^(operation_194_5523));
            operation_194_5479 <= ((operation_194_4962)^(operation_194_5486));
            operation_194_5489 <= ((operation_194_5490)^(operation_194_5494));
            operation_194_5490 <= ((operation_194_5493)^(operation_194_5524));
            operation_194_5491 <= ((operation_194_5492)^(operation_194_5498));
            operation_194_5492 <= ((operation_194_5497)^(operation_194_5528));
            operation_194_5504 <= ((operation_194_5021)^(operation_194_5519));
            operation_194_5506 <= ((operation_194_5020)^(operation_194_5517));
            operation_194_5521_latch <= (operation_194_5521);
            operation_194_5522_latch <= (operation_194_5522);
            operation_194_5531_latch <= (operation_194_5531);
            operation_194_5532_latch <= (operation_194_5532);
            operation_194_5533_latch <= (operation_194_5533);
            operation_194_5534_latch <= (operation_194_5534);
            operation_194_5535_latch <= (operation_194_5535);
            operation_194_5536_latch <= (operation_194_5536);
            operation_194_5537_latch <= (operation_194_5537);
            operation_194_5538_latch <= (operation_194_5538);
            operation_194_5539_latch <= (operation_194_5539);
            operation_194_5540_latch <= (operation_194_5540);
            operation_194_5541_latch <= (operation_194_5541);
            operation_194_5542_latch <= (operation_194_5542);
            operation_194_5543_latch <= (operation_194_5543);
            operation_194_5544_latch <= (operation_194_5544);
            operation_194_5545_latch <= (operation_194_5545);
            operation_194_5546_latch <= (operation_194_5546);
            operation_194_5547_latch <= (operation_194_5547);
            operation_194_5548_latch <= (operation_194_5548);
            operation_194_4703 <= ((operation_194_4724)^(operation_194_4704));
            operation_194_4707 <= ((operation_194_4275)^(operation_194_4731));
            operation_194_4709 <= ((operation_194_4730)^(operation_194_4863));
            operation_194_4711 <= ((operation_194_4729)^(operation_194_4962));
            operation_194_4713 <= ((operation_194_4728)^(operation_194_4803));
            operation_194_4715 <= ((operation_194_4727)^(operation_194_4862));
            operation_194_4717 <= ((operation_194_4726)^(operation_194_4731));
            operation_194_4719 <= ((operation_194_4725)^(operation_194_4802));
            operation_194_4721 <= ((operation_194_4723)^(operation_194_4722));
            operation_194_4733 <= ((operation_194_5070)^(operation_194_4781));
            operation_194_4735 <= ((operation_194_5071)^(operation_194_4780));
            operation_194_4737 <= ((operation_194_5068)^(operation_194_4779));
            operation_194_4739 <= ((operation_194_5069)^(operation_194_4778));
            operation_194_4741 <= ((operation_194_5066)^(operation_194_4777));
            operation_194_4743 <= ((operation_194_5067)^(operation_194_4776));
            operation_194_4745 <= ((operation_194_5064)^(operation_194_4775));
            operation_194_4747 <= ((operation_194_5065)^(operation_194_4774));
            operation_194_4749 <= ((operation_194_4773)^(operation_194_5021));
            operation_194_4751 <= ((operation_194_4772)^(operation_194_5020));
            operation_194_4753 <= ((operation_194_4771)^(operation_194_4901));
            operation_194_4755 <= ((operation_194_4770)^(operation_194_4900));
            operation_194_4757 <= ((operation_194_4769)^(operation_194_4833));
            operation_194_4759 <= ((operation_194_4768)^(operation_194_4832));
            operation_194_4761 <= ((operation_194_4767)^(operation_194_4766));
            operation_194_4763 <= ((operation_194_4765)^(operation_194_4764));
            operation_194_4783 <= ((operation_194_5101)^(operation_194_4811));
            operation_194_4785 <= ((operation_194_5100)^(operation_194_4810));
            operation_194_4787 <= ((operation_194_5099)^(operation_194_4809));
            operation_194_4789 <= ((operation_194_5098)^(operation_194_4808));
            operation_194_4791 <= ((operation_194_5097)^(operation_194_4807));
            operation_194_4793 <= ((operation_194_5096)^(operation_194_4806));
            operation_194_4795 <= ((operation_194_5095)^(operation_194_4805));
            operation_194_4797 <= ((operation_194_5094)^(operation_194_4804));
            operation_194_4799 <= ((operation_194_4302)^(operation_194_4803));
            operation_194_4801 <= ((operation_194_4293)^(operation_194_4802));
            operation_194_4813 <= ((operation_194_4841)^(operation_194_4965));
            operation_194_4815 <= ((operation_194_4840)^(operation_194_4965));
            operation_194_4817 <= ((operation_194_4839)^(operation_194_5024));
            operation_194_4819 <= ((operation_194_4838)^(operation_194_5024));
            operation_194_4821 <= ((operation_194_4837)^(operation_194_4964));
            operation_194_4823 <= ((operation_194_4836)^(operation_194_4964));
            operation_194_4825 <= ((operation_194_4835)^(operation_194_5023));
            operation_194_4827 <= ((operation_194_4834)^(operation_194_5023));
            operation_194_4829 <= ((operation_194_4337)^(operation_194_4833));
            operation_194_4831 <= ((operation_194_4335)^(operation_194_4832));
            operation_194_4843 <= ((operation_194_4871)^(operation_194_4965));
            operation_194_4845 <= ((operation_194_4870)^(operation_194_4965));
            operation_194_4847 <= ((operation_194_4869)^(operation_194_5024));
            operation_194_4849 <= ((operation_194_4868)^(operation_194_5024));
            operation_194_4851 <= ((operation_194_4867)^(operation_194_4964));
            operation_194_4853 <= ((operation_194_4866)^(operation_194_4964));
            operation_194_4855 <= ((operation_194_4865)^(operation_194_5023));
            operation_194_4857 <= ((operation_194_4864)^(operation_194_5023));
            operation_194_4859 <= ((operation_194_4374)^(operation_194_4863));
            operation_194_4861 <= ((operation_194_4373)^(operation_194_4862));
            operation_194_4873 <= ((operation_194_4932)^(operation_194_4874));
            operation_194_4874 <= ((operation_194_4930)*(operation_194_5597));
            operation_194_4876 <= ((operation_194_4928)^(operation_194_4877));
            operation_194_4877 <= ((operation_194_4926)*(operation_194_5597));
            operation_194_4879 <= ((operation_194_4924)^(operation_194_4880));
            operation_194_4880 <= ((operation_194_4922)*(operation_194_5597));
            operation_194_4882 <= ((operation_194_4920)^(operation_194_4883));
            operation_194_4883 <= ((operation_194_4918)*(operation_194_5597));
            operation_194_4885 <= ((operation_194_4916)^(operation_194_4886));
            operation_194_4886 <= ((operation_194_4914)*(operation_194_5597));
            operation_194_4888 <= ((operation_194_4912)^(operation_194_4889));
            operation_194_4889 <= ((operation_194_4910)*(operation_194_5597));
            operation_194_4891 <= ((operation_194_4908)^(operation_194_4892));
            operation_194_4892 <= ((operation_194_4906)*(operation_194_5597));
            operation_194_4894 <= ((operation_194_4904)^(operation_194_4895));
            operation_194_4895 <= ((operation_194_4902)*(operation_194_5597));
            operation_194_4897 <= ((operation_194_4404)^(operation_194_4901));
            operation_194_4899 <= ((operation_194_4403)^(operation_194_4900));
            operation_194_4902 <= ((operation_194_4903)&(operation_194_5557));
            operation_194_4903 <= ((operation_194_4905)>>(operation_194_2119));
            operation_194_4904 <= ((operation_194_4905)<<(operation_194_5557));
            operation_194_4906 <= ((operation_194_4907)&(operation_194_5557));
            operation_194_4907 <= ((operation_194_4909)>>(operation_194_2119));
            operation_194_4908 <= ((operation_194_4909)<<(operation_194_5557));
            operation_194_4910 <= ((operation_194_4911)&(operation_194_5557));
            operation_194_4911 <= ((operation_194_4913)>>(operation_194_2119));
            operation_194_4912 <= ((operation_194_4913)<<(operation_194_5557));
            operation_194_4914 <= ((operation_194_4915)&(operation_194_5557));
            operation_194_4915 <= ((operation_194_4917)>>(operation_194_2119));
            operation_194_4916 <= ((operation_194_4917)<<(operation_194_5557));
            operation_194_4918 <= ((operation_194_4919)&(operation_194_5557));
            operation_194_4919 <= ((operation_194_4921)>>(operation_194_2119));
            operation_194_4920 <= ((operation_194_4921)<<(operation_194_5557));
            operation_194_4922 <= ((operation_194_4923)&(operation_194_5557));
            operation_194_4923 <= ((operation_194_4925)>>(operation_194_2119));
            operation_194_4924 <= ((operation_194_4925)<<(operation_194_5557));
            operation_194_4926 <= ((operation_194_4927)&(operation_194_5557));
            operation_194_4927 <= ((operation_194_4929)>>(operation_194_2119));
            operation_194_4928 <= ((operation_194_4929)<<(operation_194_5557));
            operation_194_4930 <= ((operation_194_4931)&(operation_194_5557));
            operation_194_4931 <= ((operation_194_4933)>>(operation_194_2119));
            operation_194_4932 <= ((operation_194_4933)<<(operation_194_5557));
            operation_194_4935 <= ((operation_194_4996)^(operation_194_4936));
            operation_194_4936 <= ((operation_194_4994)*(operation_194_5597));
            operation_194_4938 <= ((operation_194_4992)^(operation_194_4939));
            operation_194_4939 <= ((operation_194_4990)*(operation_194_5597));
            operation_194_4941 <= ((operation_194_4988)^(operation_194_4942));
            operation_194_4942 <= ((operation_194_4986)*(operation_194_5597));
            operation_194_4944 <= ((operation_194_4984)^(operation_194_4945));
            operation_194_4945 <= ((operation_194_4982)*(operation_194_5597));
            operation_194_4947 <= ((operation_194_4980)^(operation_194_4948));
            operation_194_4948 <= ((operation_194_4978)*(operation_194_5597));
            operation_194_4950 <= ((operation_194_4976)^(operation_194_4951));
            operation_194_4951 <= ((operation_194_4974)*(operation_194_5597));
            operation_194_4953 <= ((operation_194_4972)^(operation_194_4954));
            operation_194_4954 <= ((operation_194_4970)*(operation_194_5597));
            operation_194_4956 <= ((operation_194_4968)^(operation_194_4957));
            operation_194_4957 <= ((operation_194_4966)*(operation_194_5597));
            operation_194_4959 <= ((operation_194_4434)^(operation_194_4963));
            operation_194_4961 <= ((operation_194_4433)^(operation_194_4962));
            operation_194_4966 <= ((operation_194_4967)&(operation_194_5557));
            operation_194_4967 <= ((operation_194_4969)>>(operation_194_2119));
            operation_194_4968 <= ((operation_194_4969)<<(operation_194_5557));
            operation_194_4970 <= ((operation_194_4971)&(operation_194_5557));
            operation_194_4971 <= ((operation_194_4973)>>(operation_194_2119));
            operation_194_4972 <= ((operation_194_4973)<<(operation_194_5557));
            operation_194_4974 <= ((operation_194_4975)&(operation_194_5557));
            operation_194_4975 <= ((operation_194_4977)>>(operation_194_2119));
            operation_194_4976 <= ((operation_194_4977)<<(operation_194_5557));
            operation_194_4978 <= ((operation_194_4979)&(operation_194_5557));
            operation_194_4979 <= ((operation_194_4981)>>(operation_194_2119));
            operation_194_4980 <= ((operation_194_4981)<<(operation_194_5557));
            operation_194_4982 <= ((operation_194_4983)&(operation_194_5557));
            operation_194_4983 <= ((operation_194_4985)>>(operation_194_2119));
            operation_194_4984 <= ((operation_194_4985)<<(operation_194_5557));
            operation_194_4986 <= ((operation_194_4987)&(operation_194_5557));
            operation_194_4987 <= ((operation_194_4989)>>(operation_194_2119));
            operation_194_4988 <= ((operation_194_4989)<<(operation_194_5557));
            operation_194_4990 <= ((operation_194_4991)&(operation_194_5557));
            operation_194_4991 <= ((operation_194_4993)>>(operation_194_2119));
            operation_194_4992 <= ((operation_194_4993)<<(operation_194_5557));
            operation_194_4994 <= ((operation_194_4995)&(operation_194_5557));
            operation_194_4995 <= ((operation_194_4997)>>(operation_194_2119));
            operation_194_4996 <= ((operation_194_4997)<<(operation_194_5557));
            operation_194_5000 <= ((operation_194_5071)^(operation_194_5100));
            operation_194_5003 <= ((operation_194_5069)^(operation_194_5098));
            operation_194_5006 <= ((operation_194_5067)^(operation_194_5096));
            operation_194_5009 <= ((operation_194_5065)^(operation_194_5094));
            operation_194_5011 <= ((operation_194_5027)^(operation_194_5100));
            operation_194_5013 <= ((operation_194_5025)^(operation_194_5096));
            operation_194_5015 <= ((operation_194_5022)^(operation_194_5592));
            operation_194_5017 <= ((operation_194_4472)^(operation_194_5021));
            operation_194_5019 <= ((operation_194_4471)^(operation_194_5020));
            operation_194_5025 <= ((operation_194_5026)^(operation_194_5067));
            operation_194_5026 <= ((operation_194_5066)^(operation_194_5097));
            operation_194_5027 <= ((operation_194_5028)^(operation_194_5071));
            operation_194_5028 <= ((operation_194_5070)^(operation_194_5101));
            operation_194_5030 <= ((operation_194_5101)^(operation_194_5071));
            operation_194_5032 <= ((operation_194_5100)^(operation_194_5070));
            operation_194_5034 <= ((operation_194_5099)^(operation_194_5069));
            operation_194_5036 <= ((operation_194_5098)^(operation_194_5068));
            operation_194_5038 <= ((operation_194_5097)^(operation_194_5067));
            operation_194_5040 <= ((operation_194_5096)^(operation_194_5066));
            operation_194_5042 <= ((operation_194_5095)^(operation_194_5065));
            operation_194_5044 <= ((operation_194_5094)^(operation_194_5064));
            operation_194_5046 <= ((operation_194_5062)^(operation_194_5098));
            operation_194_5048 <= ((operation_194_5060)^(operation_194_5094));
            operation_194_5050 <= ((operation_194_4533)^(operation_194_5057));
            operation_194_5060 <= ((operation_194_5061)^(operation_194_5065));
            operation_194_5061 <= ((operation_194_5064)^(operation_194_5095));
            operation_194_5062 <= ((operation_194_5063)^(operation_194_5069));
            operation_194_5063 <= ((operation_194_5068)^(operation_194_5099));
            operation_194_5075 <= ((operation_194_4592)^(operation_194_5090));
            operation_194_5077 <= ((operation_194_4591)^(operation_194_5088));
            operation_194_5092_latch <= (operation_194_5092);
            operation_194_5093_latch <= (operation_194_5093);
            operation_194_5102_latch <= (operation_194_5102);
            operation_194_5103_latch <= (operation_194_5103);
            operation_194_5104_latch <= (operation_194_5104);
            operation_194_5105_latch <= (operation_194_5105);
            operation_194_5106_latch <= (operation_194_5106);
            operation_194_5107_latch <= (operation_194_5107);
            operation_194_5108_latch <= (operation_194_5108);
            operation_194_5109_latch <= (operation_194_5109);
            operation_194_5110_latch <= (operation_194_5110);
            operation_194_5111_latch <= (operation_194_5111);
            operation_194_5112_latch <= (operation_194_5112);
            operation_194_5113_latch <= (operation_194_5113);
            operation_194_5114_latch <= (operation_194_5114);
            operation_194_5115_latch <= (operation_194_5115);
            operation_194_5116_latch <= (operation_194_5116);
            operation_194_5117_latch <= (operation_194_5117);
            operation_194_5118_latch <= (operation_194_5118);
            operation_194_5119_latch <= (operation_194_5119);
            operation_194_4274 <= ((operation_194_4295)^(operation_194_4275));
            operation_194_4278 <= ((operation_194_3846)^(operation_194_4302));
            operation_194_4280 <= ((operation_194_4301)^(operation_194_4434));
            operation_194_4282 <= ((operation_194_4300)^(operation_194_4533));
            operation_194_4284 <= ((operation_194_4299)^(operation_194_4374));
            operation_194_4286 <= ((operation_194_4298)^(operation_194_4433));
            operation_194_4288 <= ((operation_194_4297)^(operation_194_4302));
            operation_194_4290 <= ((operation_194_4296)^(operation_194_4373));
            operation_194_4292 <= ((operation_194_4294)^(operation_194_4293));
            operation_194_4304 <= ((operation_194_4641)^(operation_194_4352));
            operation_194_4306 <= ((operation_194_4642)^(operation_194_4351));
            operation_194_4308 <= ((operation_194_4639)^(operation_194_4350));
            operation_194_4310 <= ((operation_194_4640)^(operation_194_4349));
            operation_194_4312 <= ((operation_194_4637)^(operation_194_4348));
            operation_194_4314 <= ((operation_194_4638)^(operation_194_4347));
            operation_194_4316 <= ((operation_194_4635)^(operation_194_4346));
            operation_194_4318 <= ((operation_194_4636)^(operation_194_4345));
            operation_194_4320 <= ((operation_194_4344)^(operation_194_4592));
            operation_194_4322 <= ((operation_194_4343)^(operation_194_4591));
            operation_194_4324 <= ((operation_194_4342)^(operation_194_4472));
            operation_194_4326 <= ((operation_194_4341)^(operation_194_4471));
            operation_194_4328 <= ((operation_194_4340)^(operation_194_4404));
            operation_194_4330 <= ((operation_194_4339)^(operation_194_4403));
            operation_194_4332 <= ((operation_194_4338)^(operation_194_4337));
            operation_194_4334 <= ((operation_194_4336)^(operation_194_4335));
            operation_194_4354 <= ((operation_194_4672)^(operation_194_4382));
            operation_194_4356 <= ((operation_194_4671)^(operation_194_4381));
            operation_194_4358 <= ((operation_194_4670)^(operation_194_4380));
            operation_194_4360 <= ((operation_194_4669)^(operation_194_4379));
            operation_194_4362 <= ((operation_194_4668)^(operation_194_4378));
            operation_194_4364 <= ((operation_194_4667)^(operation_194_4377));
            operation_194_4366 <= ((operation_194_4666)^(operation_194_4376));
            operation_194_4368 <= ((operation_194_4665)^(operation_194_4375));
            operation_194_4370 <= ((operation_194_3873)^(operation_194_4374));
            operation_194_4372 <= ((operation_194_3864)^(operation_194_4373));
            operation_194_4384 <= ((operation_194_4412)^(operation_194_4536));
            operation_194_4386 <= ((operation_194_4411)^(operation_194_4536));
            operation_194_4388 <= ((operation_194_4410)^(operation_194_4595));
            operation_194_4390 <= ((operation_194_4409)^(operation_194_4595));
            operation_194_4392 <= ((operation_194_4408)^(operation_194_4535));
            operation_194_4394 <= ((operation_194_4407)^(operation_194_4535));
            operation_194_4396 <= ((operation_194_4406)^(operation_194_4594));
            operation_194_4398 <= ((operation_194_4405)^(operation_194_4594));
            operation_194_4400 <= ((operation_194_3908)^(operation_194_4404));
            operation_194_4402 <= ((operation_194_3906)^(operation_194_4403));
            operation_194_4414 <= ((operation_194_4442)^(operation_194_4536));
            operation_194_4416 <= ((operation_194_4441)^(operation_194_4536));
            operation_194_4418 <= ((operation_194_4440)^(operation_194_4595));
            operation_194_4420 <= ((operation_194_4439)^(operation_194_4595));
            operation_194_4422 <= ((operation_194_4438)^(operation_194_4535));
            operation_194_4424 <= ((operation_194_4437)^(operation_194_4535));
            operation_194_4426 <= ((operation_194_4436)^(operation_194_4594));
            operation_194_4428 <= ((operation_194_4435)^(operation_194_4594));
            operation_194_4430 <= ((operation_194_3945)^(operation_194_4434));
            operation_194_4432 <= ((operation_194_3944)^(operation_194_4433));
            operation_194_4444 <= ((operation_194_4503)^(operation_194_4445));
            operation_194_4445 <= ((operation_194_4501)*(operation_194_5597));
            operation_194_4447 <= ((operation_194_4499)^(operation_194_4448));
            operation_194_4448 <= ((operation_194_4497)*(operation_194_5597));
            operation_194_4450 <= ((operation_194_4495)^(operation_194_4451));
            operation_194_4451 <= ((operation_194_4493)*(operation_194_5597));
            operation_194_4453 <= ((operation_194_4491)^(operation_194_4454));
            operation_194_4454 <= ((operation_194_4489)*(operation_194_5597));
            operation_194_4456 <= ((operation_194_4487)^(operation_194_4457));
            operation_194_4457 <= ((operation_194_4485)*(operation_194_5597));
            operation_194_4459 <= ((operation_194_4483)^(operation_194_4460));
            operation_194_4460 <= ((operation_194_4481)*(operation_194_5597));
            operation_194_4462 <= ((operation_194_4479)^(operation_194_4463));
            operation_194_4463 <= ((operation_194_4477)*(operation_194_5597));
            operation_194_4465 <= ((operation_194_4475)^(operation_194_4466));
            operation_194_4466 <= ((operation_194_4473)*(operation_194_5597));
            operation_194_4468 <= ((operation_194_3975)^(operation_194_4472));
            operation_194_4470 <= ((operation_194_3974)^(operation_194_4471));
            operation_194_4473 <= ((operation_194_4474)&(operation_194_5557));
            operation_194_4474 <= ((operation_194_4476)>>(operation_194_2119));
            operation_194_4475 <= ((operation_194_4476)<<(operation_194_5557));
            operation_194_4477 <= ((operation_194_4478)&(operation_194_5557));
            operation_194_4478 <= ((operation_194_4480)>>(operation_194_2119));
            operation_194_4479 <= ((operation_194_4480)<<(operation_194_5557));
            operation_194_4481 <= ((operation_194_4482)&(operation_194_5557));
            operation_194_4482 <= ((operation_194_4484)>>(operation_194_2119));
            operation_194_4483 <= ((operation_194_4484)<<(operation_194_5557));
            operation_194_4485 <= ((operation_194_4486)&(operation_194_5557));
            operation_194_4486 <= ((operation_194_4488)>>(operation_194_2119));
            operation_194_4487 <= ((operation_194_4488)<<(operation_194_5557));
            operation_194_4489 <= ((operation_194_4490)&(operation_194_5557));
            operation_194_4490 <= ((operation_194_4492)>>(operation_194_2119));
            operation_194_4491 <= ((operation_194_4492)<<(operation_194_5557));
            operation_194_4493 <= ((operation_194_4494)&(operation_194_5557));
            operation_194_4494 <= ((operation_194_4496)>>(operation_194_2119));
            operation_194_4495 <= ((operation_194_4496)<<(operation_194_5557));
            operation_194_4497 <= ((operation_194_4498)&(operation_194_5557));
            operation_194_4498 <= ((operation_194_4500)>>(operation_194_2119));
            operation_194_4499 <= ((operation_194_4500)<<(operation_194_5557));
            operation_194_4501 <= ((operation_194_4502)&(operation_194_5557));
            operation_194_4502 <= ((operation_194_4504)>>(operation_194_2119));
            operation_194_4503 <= ((operation_194_4504)<<(operation_194_5557));
            operation_194_4506 <= ((operation_194_4567)^(operation_194_4507));
            operation_194_4507 <= ((operation_194_4565)*(operation_194_5597));
            operation_194_4509 <= ((operation_194_4563)^(operation_194_4510));
            operation_194_4510 <= ((operation_194_4561)*(operation_194_5597));
            operation_194_4512 <= ((operation_194_4559)^(operation_194_4513));
            operation_194_4513 <= ((operation_194_4557)*(operation_194_5597));
            operation_194_4515 <= ((operation_194_4555)^(operation_194_4516));
            operation_194_4516 <= ((operation_194_4553)*(operation_194_5597));
            operation_194_4518 <= ((operation_194_4551)^(operation_194_4519));
            operation_194_4519 <= ((operation_194_4549)*(operation_194_5597));
            operation_194_4521 <= ((operation_194_4547)^(operation_194_4522));
            operation_194_4522 <= ((operation_194_4545)*(operation_194_5597));
            operation_194_4524 <= ((operation_194_4543)^(operation_194_4525));
            operation_194_4525 <= ((operation_194_4541)*(operation_194_5597));
            operation_194_4527 <= ((operation_194_4539)^(operation_194_4528));
            operation_194_4528 <= ((operation_194_4537)*(operation_194_5597));
            operation_194_4530 <= ((operation_194_4005)^(operation_194_4534));
            operation_194_4532 <= ((operation_194_4004)^(operation_194_4533));
            operation_194_4537 <= ((operation_194_4538)&(operation_194_5557));
            operation_194_4538 <= ((operation_194_4540)>>(operation_194_2119));
            operation_194_4539 <= ((operation_194_4540)<<(operation_194_5557));
            operation_194_4541 <= ((operation_194_4542)&(operation_194_5557));
            operation_194_4542 <= ((operation_194_4544)>>(operation_194_2119));
            operation_194_4543 <= ((operation_194_4544)<<(operation_194_5557));
            operation_194_4545 <= ((operation_194_4546)&(operation_194_5557));
            operation_194_4546 <= ((operation_194_4548)>>(operation_194_2119));
            operation_194_4547 <= ((operation_194_4548)<<(operation_194_5557));
            operation_194_4549 <= ((operation_194_4550)&(operation_194_5557));
            operation_194_4550 <= ((operation_194_4552)>>(operation_194_2119));
            operation_194_4551 <= ((operation_194_4552)<<(operation_194_5557));
            operation_194_4553 <= ((operation_194_4554)&(operation_194_5557));
            operation_194_4554 <= ((operation_194_4556)>>(operation_194_2119));
            operation_194_4555 <= ((operation_194_4556)<<(operation_194_5557));
            operation_194_4557 <= ((operation_194_4558)&(operation_194_5557));
            operation_194_4558 <= ((operation_194_4560)>>(operation_194_2119));
            operation_194_4559 <= ((operation_194_4560)<<(operation_194_5557));
            operation_194_4561 <= ((operation_194_4562)&(operation_194_5557));
            operation_194_4562 <= ((operation_194_4564)>>(operation_194_2119));
            operation_194_4563 <= ((operation_194_4564)<<(operation_194_5557));
            operation_194_4565 <= ((operation_194_4566)&(operation_194_5557));
            operation_194_4566 <= ((operation_194_4568)>>(operation_194_2119));
            operation_194_4567 <= ((operation_194_4568)<<(operation_194_5557));
            operation_194_4571 <= ((operation_194_4642)^(operation_194_4671));
            operation_194_4574 <= ((operation_194_4640)^(operation_194_4669));
            operation_194_4577 <= ((operation_194_4638)^(operation_194_4667));
            operation_194_4580 <= ((operation_194_4636)^(operation_194_4665));
            operation_194_4582 <= ((operation_194_4598)^(operation_194_4671));
            operation_194_4584 <= ((operation_194_4596)^(operation_194_4667));
            operation_194_4586 <= ((operation_194_4593)^(operation_194_5587));
            operation_194_4588 <= ((operation_194_4043)^(operation_194_4592));
            operation_194_4590 <= ((operation_194_4042)^(operation_194_4591));
            operation_194_4596 <= ((operation_194_4597)^(operation_194_4638));
            operation_194_4597 <= ((operation_194_4637)^(operation_194_4668));
            operation_194_4598 <= ((operation_194_4599)^(operation_194_4642));
            operation_194_4599 <= ((operation_194_4641)^(operation_194_4672));
            operation_194_4601 <= ((operation_194_4672)^(operation_194_4642));
            operation_194_4603 <= ((operation_194_4671)^(operation_194_4641));
            operation_194_4605 <= ((operation_194_4670)^(operation_194_4640));
            operation_194_4607 <= ((operation_194_4669)^(operation_194_4639));
            operation_194_4609 <= ((operation_194_4668)^(operation_194_4638));
            operation_194_4611 <= ((operation_194_4667)^(operation_194_4637));
            operation_194_4613 <= ((operation_194_4666)^(operation_194_4636));
            operation_194_4615 <= ((operation_194_4665)^(operation_194_4635));
            operation_194_4617 <= ((operation_194_4633)^(operation_194_4669));
            operation_194_4619 <= ((operation_194_4631)^(operation_194_4665));
            operation_194_4621 <= ((operation_194_4104)^(operation_194_4628));
            operation_194_4631 <= ((operation_194_4632)^(operation_194_4636));
            operation_194_4632 <= ((operation_194_4635)^(operation_194_4666));
            operation_194_4633 <= ((operation_194_4634)^(operation_194_4640));
            operation_194_4634 <= ((operation_194_4639)^(operation_194_4670));
            operation_194_4646 <= ((operation_194_4163)^(operation_194_4661));
            operation_194_4648 <= ((operation_194_4162)^(operation_194_4659));
            operation_194_4663_latch <= (operation_194_4663);
            operation_194_4664_latch <= (operation_194_4664);
            operation_194_4673_latch <= (operation_194_4673);
            operation_194_4674_latch <= (operation_194_4674);
            operation_194_4675_latch <= (operation_194_4675);
            operation_194_4676_latch <= (operation_194_4676);
            operation_194_4677_latch <= (operation_194_4677);
            operation_194_4678_latch <= (operation_194_4678);
            operation_194_4679_latch <= (operation_194_4679);
            operation_194_4680_latch <= (operation_194_4680);
            operation_194_4681_latch <= (operation_194_4681);
            operation_194_4682_latch <= (operation_194_4682);
            operation_194_4683_latch <= (operation_194_4683);
            operation_194_4684_latch <= (operation_194_4684);
            operation_194_4685_latch <= (operation_194_4685);
            operation_194_4686_latch <= (operation_194_4686);
            operation_194_4687_latch <= (operation_194_4687);
            operation_194_4688_latch <= (operation_194_4688);
            operation_194_4689_latch <= (operation_194_4689);
            operation_194_4690_latch <= (operation_194_4690);
            operation_194_3845 <= ((operation_194_3866)^(operation_194_3846));
            operation_194_3849 <= ((operation_194_3417)^(operation_194_3873));
            operation_194_3851 <= ((operation_194_3872)^(operation_194_4005));
            operation_194_3853 <= ((operation_194_3871)^(operation_194_4104));
            operation_194_3855 <= ((operation_194_3870)^(operation_194_3945));
            operation_194_3857 <= ((operation_194_3869)^(operation_194_4004));
            operation_194_3859 <= ((operation_194_3868)^(operation_194_3873));
            operation_194_3861 <= ((operation_194_3867)^(operation_194_3944));
            operation_194_3863 <= ((operation_194_3865)^(operation_194_3864));
            operation_194_3875 <= ((operation_194_4212)^(operation_194_3923));
            operation_194_3877 <= ((operation_194_4213)^(operation_194_3922));
            operation_194_3879 <= ((operation_194_4210)^(operation_194_3921));
            operation_194_3881 <= ((operation_194_4211)^(operation_194_3920));
            operation_194_3883 <= ((operation_194_4208)^(operation_194_3919));
            operation_194_3885 <= ((operation_194_4209)^(operation_194_3918));
            operation_194_3887 <= ((operation_194_4206)^(operation_194_3917));
            operation_194_3889 <= ((operation_194_4207)^(operation_194_3916));
            operation_194_3891 <= ((operation_194_3915)^(operation_194_4163));
            operation_194_3893 <= ((operation_194_3914)^(operation_194_4162));
            operation_194_3895 <= ((operation_194_3913)^(operation_194_4043));
            operation_194_3897 <= ((operation_194_3912)^(operation_194_4042));
            operation_194_3899 <= ((operation_194_3911)^(operation_194_3975));
            operation_194_3901 <= ((operation_194_3910)^(operation_194_3974));
            operation_194_3903 <= ((operation_194_3909)^(operation_194_3908));
            operation_194_3905 <= ((operation_194_3907)^(operation_194_3906));
            operation_194_3925 <= ((operation_194_4243)^(operation_194_3953));
            operation_194_3927 <= ((operation_194_4242)^(operation_194_3952));
            operation_194_3929 <= ((operation_194_4241)^(operation_194_3951));
            operation_194_3931 <= ((operation_194_4240)^(operation_194_3950));
            operation_194_3933 <= ((operation_194_4239)^(operation_194_3949));
            operation_194_3935 <= ((operation_194_4238)^(operation_194_3948));
            operation_194_3937 <= ((operation_194_4237)^(operation_194_3947));
            operation_194_3939 <= ((operation_194_4236)^(operation_194_3946));
            operation_194_3941 <= ((operation_194_3444)^(operation_194_3945));
            operation_194_3943 <= ((operation_194_3435)^(operation_194_3944));
            operation_194_3955 <= ((operation_194_3983)^(operation_194_4107));
            operation_194_3957 <= ((operation_194_3982)^(operation_194_4107));
            operation_194_3959 <= ((operation_194_3981)^(operation_194_4166));
            operation_194_3961 <= ((operation_194_3980)^(operation_194_4166));
            operation_194_3963 <= ((operation_194_3979)^(operation_194_4106));
            operation_194_3965 <= ((operation_194_3978)^(operation_194_4106));
            operation_194_3967 <= ((operation_194_3977)^(operation_194_4165));
            operation_194_3969 <= ((operation_194_3976)^(operation_194_4165));
            operation_194_3971 <= ((operation_194_3479)^(operation_194_3975));
            operation_194_3973 <= ((operation_194_3477)^(operation_194_3974));
            operation_194_3985 <= ((operation_194_4013)^(operation_194_4107));
            operation_194_3987 <= ((operation_194_4012)^(operation_194_4107));
            operation_194_3989 <= ((operation_194_4011)^(operation_194_4166));
            operation_194_3991 <= ((operation_194_4010)^(operation_194_4166));
            operation_194_3993 <= ((operation_194_4009)^(operation_194_4106));
            operation_194_3995 <= ((operation_194_4008)^(operation_194_4106));
            operation_194_3997 <= ((operation_194_4007)^(operation_194_4165));
            operation_194_3999 <= ((operation_194_4006)^(operation_194_4165));
            operation_194_4001 <= ((operation_194_3516)^(operation_194_4005));
            operation_194_4003 <= ((operation_194_3515)^(operation_194_4004));
            operation_194_4015 <= ((operation_194_4074)^(operation_194_4016));
            operation_194_4016 <= ((operation_194_4072)*(operation_194_5597));
            operation_194_4018 <= ((operation_194_4070)^(operation_194_4019));
            operation_194_4019 <= ((operation_194_4068)*(operation_194_5597));
            operation_194_4021 <= ((operation_194_4066)^(operation_194_4022));
            operation_194_4022 <= ((operation_194_4064)*(operation_194_5597));
            operation_194_4024 <= ((operation_194_4062)^(operation_194_4025));
            operation_194_4025 <= ((operation_194_4060)*(operation_194_5597));
            operation_194_4027 <= ((operation_194_4058)^(operation_194_4028));
            operation_194_4028 <= ((operation_194_4056)*(operation_194_5597));
            operation_194_4030 <= ((operation_194_4054)^(operation_194_4031));
            operation_194_4031 <= ((operation_194_4052)*(operation_194_5597));
            operation_194_4033 <= ((operation_194_4050)^(operation_194_4034));
            operation_194_4034 <= ((operation_194_4048)*(operation_194_5597));
            operation_194_4036 <= ((operation_194_4046)^(operation_194_4037));
            operation_194_4037 <= ((operation_194_4044)*(operation_194_5597));
            operation_194_4039 <= ((operation_194_3546)^(operation_194_4043));
            operation_194_4041 <= ((operation_194_3545)^(operation_194_4042));
            operation_194_4044 <= ((operation_194_4045)&(operation_194_5557));
            operation_194_4045 <= ((operation_194_4047)>>(operation_194_2119));
            operation_194_4046 <= ((operation_194_4047)<<(operation_194_5557));
            operation_194_4048 <= ((operation_194_4049)&(operation_194_5557));
            operation_194_4049 <= ((operation_194_4051)>>(operation_194_2119));
            operation_194_4050 <= ((operation_194_4051)<<(operation_194_5557));
            operation_194_4052 <= ((operation_194_4053)&(operation_194_5557));
            operation_194_4053 <= ((operation_194_4055)>>(operation_194_2119));
            operation_194_4054 <= ((operation_194_4055)<<(operation_194_5557));
            operation_194_4056 <= ((operation_194_4057)&(operation_194_5557));
            operation_194_4057 <= ((operation_194_4059)>>(operation_194_2119));
            operation_194_4058 <= ((operation_194_4059)<<(operation_194_5557));
            operation_194_4060 <= ((operation_194_4061)&(operation_194_5557));
            operation_194_4061 <= ((operation_194_4063)>>(operation_194_2119));
            operation_194_4062 <= ((operation_194_4063)<<(operation_194_5557));
            operation_194_4064 <= ((operation_194_4065)&(operation_194_5557));
            operation_194_4065 <= ((operation_194_4067)>>(operation_194_2119));
            operation_194_4066 <= ((operation_194_4067)<<(operation_194_5557));
            operation_194_4068 <= ((operation_194_4069)&(operation_194_5557));
            operation_194_4069 <= ((operation_194_4071)>>(operation_194_2119));
            operation_194_4070 <= ((operation_194_4071)<<(operation_194_5557));
            operation_194_4072 <= ((operation_194_4073)&(operation_194_5557));
            operation_194_4073 <= ((operation_194_4075)>>(operation_194_2119));
            operation_194_4074 <= ((operation_194_4075)<<(operation_194_5557));
            operation_194_4077 <= ((operation_194_4138)^(operation_194_4078));
            operation_194_4078 <= ((operation_194_4136)*(operation_194_5597));
            operation_194_4080 <= ((operation_194_4134)^(operation_194_4081));
            operation_194_4081 <= ((operation_194_4132)*(operation_194_5597));
            operation_194_4083 <= ((operation_194_4130)^(operation_194_4084));
            operation_194_4084 <= ((operation_194_4128)*(operation_194_5597));
            operation_194_4086 <= ((operation_194_4126)^(operation_194_4087));
            operation_194_4087 <= ((operation_194_4124)*(operation_194_5597));
            operation_194_4089 <= ((operation_194_4122)^(operation_194_4090));
            operation_194_4090 <= ((operation_194_4120)*(operation_194_5597));
            operation_194_4092 <= ((operation_194_4118)^(operation_194_4093));
            operation_194_4093 <= ((operation_194_4116)*(operation_194_5597));
            operation_194_4095 <= ((operation_194_4114)^(operation_194_4096));
            operation_194_4096 <= ((operation_194_4112)*(operation_194_5597));
            operation_194_4098 <= ((operation_194_4110)^(operation_194_4099));
            operation_194_4099 <= ((operation_194_4108)*(operation_194_5597));
            operation_194_4101 <= ((operation_194_3576)^(operation_194_4105));
            operation_194_4103 <= ((operation_194_3575)^(operation_194_4104));
            operation_194_4108 <= ((operation_194_4109)&(operation_194_5557));
            operation_194_4109 <= ((operation_194_4111)>>(operation_194_2119));
            operation_194_4110 <= ((operation_194_4111)<<(operation_194_5557));
            operation_194_4112 <= ((operation_194_4113)&(operation_194_5557));
            operation_194_4113 <= ((operation_194_4115)>>(operation_194_2119));
            operation_194_4114 <= ((operation_194_4115)<<(operation_194_5557));
            operation_194_4116 <= ((operation_194_4117)&(operation_194_5557));
            operation_194_4117 <= ((operation_194_4119)>>(operation_194_2119));
            operation_194_4118 <= ((operation_194_4119)<<(operation_194_5557));
            operation_194_4120 <= ((operation_194_4121)&(operation_194_5557));
            operation_194_4121 <= ((operation_194_4123)>>(operation_194_2119));
            operation_194_4122 <= ((operation_194_4123)<<(operation_194_5557));
            operation_194_4124 <= ((operation_194_4125)&(operation_194_5557));
            operation_194_4125 <= ((operation_194_4127)>>(operation_194_2119));
            operation_194_4126 <= ((operation_194_4127)<<(operation_194_5557));
            operation_194_4128 <= ((operation_194_4129)&(operation_194_5557));
            operation_194_4129 <= ((operation_194_4131)>>(operation_194_2119));
            operation_194_4130 <= ((operation_194_4131)<<(operation_194_5557));
            operation_194_4132 <= ((operation_194_4133)&(operation_194_5557));
            operation_194_4133 <= ((operation_194_4135)>>(operation_194_2119));
            operation_194_4134 <= ((operation_194_4135)<<(operation_194_5557));
            operation_194_4136 <= ((operation_194_4137)&(operation_194_5557));
            operation_194_4137 <= ((operation_194_4139)>>(operation_194_2119));
            operation_194_4138 <= ((operation_194_4139)<<(operation_194_5557));
            operation_194_4142 <= ((operation_194_4213)^(operation_194_4242));
            operation_194_4145 <= ((operation_194_4211)^(operation_194_4240));
            operation_194_4148 <= ((operation_194_4209)^(operation_194_4238));
            operation_194_4151 <= ((operation_194_4207)^(operation_194_4236));
            operation_194_4153 <= ((operation_194_4169)^(operation_194_4242));
            operation_194_4155 <= ((operation_194_4167)^(operation_194_4238));
            operation_194_4157 <= ((operation_194_4164)^(operation_194_5582));
            operation_194_4159 <= ((operation_194_3614)^(operation_194_4163));
            operation_194_4161 <= ((operation_194_3613)^(operation_194_4162));
            operation_194_4167 <= ((operation_194_4168)^(operation_194_4209));
            operation_194_4168 <= ((operation_194_4208)^(operation_194_4239));
            operation_194_4169 <= ((operation_194_4170)^(operation_194_4213));
            operation_194_4170 <= ((operation_194_4212)^(operation_194_4243));
            operation_194_4172 <= ((operation_194_4243)^(operation_194_4213));
            operation_194_4174 <= ((operation_194_4242)^(operation_194_4212));
            operation_194_4176 <= ((operation_194_4241)^(operation_194_4211));
            operation_194_4178 <= ((operation_194_4240)^(operation_194_4210));
            operation_194_4180 <= ((operation_194_4239)^(operation_194_4209));
            operation_194_4182 <= ((operation_194_4238)^(operation_194_4208));
            operation_194_4184 <= ((operation_194_4237)^(operation_194_4207));
            operation_194_4186 <= ((operation_194_4236)^(operation_194_4206));
            operation_194_4188 <= ((operation_194_4204)^(operation_194_4240));
            operation_194_4190 <= ((operation_194_4202)^(operation_194_4236));
            operation_194_4192 <= ((operation_194_3675)^(operation_194_4199));
            operation_194_4202 <= ((operation_194_4203)^(operation_194_4207));
            operation_194_4203 <= ((operation_194_4206)^(operation_194_4237));
            operation_194_4204 <= ((operation_194_4205)^(operation_194_4211));
            operation_194_4205 <= ((operation_194_4210)^(operation_194_4241));
            operation_194_4217 <= ((operation_194_3734)^(operation_194_4232));
            operation_194_4219 <= ((operation_194_3733)^(operation_194_4230));
            operation_194_4234_latch <= (operation_194_4234);
            operation_194_4235_latch <= (operation_194_4235);
            operation_194_4244_latch <= (operation_194_4244);
            operation_194_4245_latch <= (operation_194_4245);
            operation_194_4246_latch <= (operation_194_4246);
            operation_194_4247_latch <= (operation_194_4247);
            operation_194_4248_latch <= (operation_194_4248);
            operation_194_4249_latch <= (operation_194_4249);
            operation_194_4250_latch <= (operation_194_4250);
            operation_194_4251_latch <= (operation_194_4251);
            operation_194_4252_latch <= (operation_194_4252);
            operation_194_4253_latch <= (operation_194_4253);
            operation_194_4254_latch <= (operation_194_4254);
            operation_194_4255_latch <= (operation_194_4255);
            operation_194_4256_latch <= (operation_194_4256);
            operation_194_4257_latch <= (operation_194_4257);
            operation_194_4258_latch <= (operation_194_4258);
            operation_194_4259_latch <= (operation_194_4259);
            operation_194_4260_latch <= (operation_194_4260);
            operation_194_4261_latch <= (operation_194_4261);
            operation_194_3416 <= ((operation_194_3437)^(operation_194_3417));
            operation_194_3420 <= ((operation_194_2988)^(operation_194_3444));
            operation_194_3422 <= ((operation_194_3443)^(operation_194_3576));
            operation_194_3424 <= ((operation_194_3442)^(operation_194_3675));
            operation_194_3426 <= ((operation_194_3441)^(operation_194_3516));
            operation_194_3428 <= ((operation_194_3440)^(operation_194_3575));
            operation_194_3430 <= ((operation_194_3439)^(operation_194_3444));
            operation_194_3432 <= ((operation_194_3438)^(operation_194_3515));
            operation_194_3434 <= ((operation_194_3436)^(operation_194_3435));
            operation_194_3446 <= ((operation_194_3783)^(operation_194_3494));
            operation_194_3448 <= ((operation_194_3784)^(operation_194_3493));
            operation_194_3450 <= ((operation_194_3781)^(operation_194_3492));
            operation_194_3452 <= ((operation_194_3782)^(operation_194_3491));
            operation_194_3454 <= ((operation_194_3779)^(operation_194_3490));
            operation_194_3456 <= ((operation_194_3780)^(operation_194_3489));
            operation_194_3458 <= ((operation_194_3777)^(operation_194_3488));
            operation_194_3460 <= ((operation_194_3778)^(operation_194_3487));
            operation_194_3462 <= ((operation_194_3486)^(operation_194_3734));
            operation_194_3464 <= ((operation_194_3485)^(operation_194_3733));
            operation_194_3466 <= ((operation_194_3484)^(operation_194_3614));
            operation_194_3468 <= ((operation_194_3483)^(operation_194_3613));
            operation_194_3470 <= ((operation_194_3482)^(operation_194_3546));
            operation_194_3472 <= ((operation_194_3481)^(operation_194_3545));
            operation_194_3474 <= ((operation_194_3480)^(operation_194_3479));
            operation_194_3476 <= ((operation_194_3478)^(operation_194_3477));
            operation_194_3496 <= ((operation_194_3814)^(operation_194_3524));
            operation_194_3498 <= ((operation_194_3813)^(operation_194_3523));
            operation_194_3500 <= ((operation_194_3812)^(operation_194_3522));
            operation_194_3502 <= ((operation_194_3811)^(operation_194_3521));
            operation_194_3504 <= ((operation_194_3810)^(operation_194_3520));
            operation_194_3506 <= ((operation_194_3809)^(operation_194_3519));
            operation_194_3508 <= ((operation_194_3808)^(operation_194_3518));
            operation_194_3510 <= ((operation_194_3807)^(operation_194_3517));
            operation_194_3512 <= ((operation_194_3015)^(operation_194_3516));
            operation_194_3514 <= ((operation_194_3006)^(operation_194_3515));
            operation_194_3526 <= ((operation_194_3554)^(operation_194_3678));
            operation_194_3528 <= ((operation_194_3553)^(operation_194_3678));
            operation_194_3530 <= ((operation_194_3552)^(operation_194_3737));
            operation_194_3532 <= ((operation_194_3551)^(operation_194_3737));
            operation_194_3534 <= ((operation_194_3550)^(operation_194_3677));
            operation_194_3536 <= ((operation_194_3549)^(operation_194_3677));
            operation_194_3538 <= ((operation_194_3548)^(operation_194_3736));
            operation_194_3540 <= ((operation_194_3547)^(operation_194_3736));
            operation_194_3542 <= ((operation_194_3050)^(operation_194_3546));
            operation_194_3544 <= ((operation_194_3048)^(operation_194_3545));
            operation_194_3556 <= ((operation_194_3584)^(operation_194_3678));
            operation_194_3558 <= ((operation_194_3583)^(operation_194_3678));
            operation_194_3560 <= ((operation_194_3582)^(operation_194_3737));
            operation_194_3562 <= ((operation_194_3581)^(operation_194_3737));
            operation_194_3564 <= ((operation_194_3580)^(operation_194_3677));
            operation_194_3566 <= ((operation_194_3579)^(operation_194_3677));
            operation_194_3568 <= ((operation_194_3578)^(operation_194_3736));
            operation_194_3570 <= ((operation_194_3577)^(operation_194_3736));
            operation_194_3572 <= ((operation_194_3087)^(operation_194_3576));
            operation_194_3574 <= ((operation_194_3086)^(operation_194_3575));
            operation_194_3586 <= ((operation_194_3645)^(operation_194_3587));
            operation_194_3587 <= ((operation_194_3643)*(operation_194_5597));
            operation_194_3589 <= ((operation_194_3641)^(operation_194_3590));
            operation_194_3590 <= ((operation_194_3639)*(operation_194_5597));
            operation_194_3592 <= ((operation_194_3637)^(operation_194_3593));
            operation_194_3593 <= ((operation_194_3635)*(operation_194_5597));
            operation_194_3595 <= ((operation_194_3633)^(operation_194_3596));
            operation_194_3596 <= ((operation_194_3631)*(operation_194_5597));
            operation_194_3598 <= ((operation_194_3629)^(operation_194_3599));
            operation_194_3599 <= ((operation_194_3627)*(operation_194_5597));
            operation_194_3601 <= ((operation_194_3625)^(operation_194_3602));
            operation_194_3602 <= ((operation_194_3623)*(operation_194_5597));
            operation_194_3604 <= ((operation_194_3621)^(operation_194_3605));
            operation_194_3605 <= ((operation_194_3619)*(operation_194_5597));
            operation_194_3607 <= ((operation_194_3617)^(operation_194_3608));
            operation_194_3608 <= ((operation_194_3615)*(operation_194_5597));
            operation_194_3610 <= ((operation_194_3117)^(operation_194_3614));
            operation_194_3612 <= ((operation_194_3116)^(operation_194_3613));
            operation_194_3615 <= ((operation_194_3616)&(operation_194_5557));
            operation_194_3616 <= ((operation_194_3618)>>(operation_194_2119));
            operation_194_3617 <= ((operation_194_3618)<<(operation_194_5557));
            operation_194_3619 <= ((operation_194_3620)&(operation_194_5557));
            operation_194_3620 <= ((operation_194_3622)>>(operation_194_2119));
            operation_194_3621 <= ((operation_194_3622)<<(operation_194_5557));
            operation_194_3623 <= ((operation_194_3624)&(operation_194_5557));
            operation_194_3624 <= ((operation_194_3626)>>(operation_194_2119));
            operation_194_3625 <= ((operation_194_3626)<<(operation_194_5557));
            operation_194_3627 <= ((operation_194_3628)&(operation_194_5557));
            operation_194_3628 <= ((operation_194_3630)>>(operation_194_2119));
            operation_194_3629 <= ((operation_194_3630)<<(operation_194_5557));
            operation_194_3631 <= ((operation_194_3632)&(operation_194_5557));
            operation_194_3632 <= ((operation_194_3634)>>(operation_194_2119));
            operation_194_3633 <= ((operation_194_3634)<<(operation_194_5557));
            operation_194_3635 <= ((operation_194_3636)&(operation_194_5557));
            operation_194_3636 <= ((operation_194_3638)>>(operation_194_2119));
            operation_194_3637 <= ((operation_194_3638)<<(operation_194_5557));
            operation_194_3639 <= ((operation_194_3640)&(operation_194_5557));
            operation_194_3640 <= ((operation_194_3642)>>(operation_194_2119));
            operation_194_3641 <= ((operation_194_3642)<<(operation_194_5557));
            operation_194_3643 <= ((operation_194_3644)&(operation_194_5557));
            operation_194_3644 <= ((operation_194_3646)>>(operation_194_2119));
            operation_194_3645 <= ((operation_194_3646)<<(operation_194_5557));
            operation_194_3648 <= ((operation_194_3709)^(operation_194_3649));
            operation_194_3649 <= ((operation_194_3707)*(operation_194_5597));
            operation_194_3651 <= ((operation_194_3705)^(operation_194_3652));
            operation_194_3652 <= ((operation_194_3703)*(operation_194_5597));
            operation_194_3654 <= ((operation_194_3701)^(operation_194_3655));
            operation_194_3655 <= ((operation_194_3699)*(operation_194_5597));
            operation_194_3657 <= ((operation_194_3697)^(operation_194_3658));
            operation_194_3658 <= ((operation_194_3695)*(operation_194_5597));
            operation_194_3660 <= ((operation_194_3693)^(operation_194_3661));
            operation_194_3661 <= ((operation_194_3691)*(operation_194_5597));
            operation_194_3663 <= ((operation_194_3689)^(operation_194_3664));
            operation_194_3664 <= ((operation_194_3687)*(operation_194_5597));
            operation_194_3666 <= ((operation_194_3685)^(operation_194_3667));
            operation_194_3667 <= ((operation_194_3683)*(operation_194_5597));
            operation_194_3669 <= ((operation_194_3681)^(operation_194_3670));
            operation_194_3670 <= ((operation_194_3679)*(operation_194_5597));
            operation_194_3672 <= ((operation_194_3147)^(operation_194_3676));
            operation_194_3674 <= ((operation_194_3146)^(operation_194_3675));
            operation_194_3679 <= ((operation_194_3680)&(operation_194_5557));
            operation_194_3680 <= ((operation_194_3682)>>(operation_194_2119));
            operation_194_3681 <= ((operation_194_3682)<<(operation_194_5557));
            operation_194_3683 <= ((operation_194_3684)&(operation_194_5557));
            operation_194_3684 <= ((operation_194_3686)>>(operation_194_2119));
            operation_194_3685 <= ((operation_194_3686)<<(operation_194_5557));
            operation_194_3687 <= ((operation_194_3688)&(operation_194_5557));
            operation_194_3688 <= ((operation_194_3690)>>(operation_194_2119));
            operation_194_3689 <= ((operation_194_3690)<<(operation_194_5557));
            operation_194_3691 <= ((operation_194_3692)&(operation_194_5557));
            operation_194_3692 <= ((operation_194_3694)>>(operation_194_2119));
            operation_194_3693 <= ((operation_194_3694)<<(operation_194_5557));
            operation_194_3695 <= ((operation_194_3696)&(operation_194_5557));
            operation_194_3696 <= ((operation_194_3698)>>(operation_194_2119));
            operation_194_3697 <= ((operation_194_3698)<<(operation_194_5557));
            operation_194_3699 <= ((operation_194_3700)&(operation_194_5557));
            operation_194_3700 <= ((operation_194_3702)>>(operation_194_2119));
            operation_194_3701 <= ((operation_194_3702)<<(operation_194_5557));
            operation_194_3703 <= ((operation_194_3704)&(operation_194_5557));
            operation_194_3704 <= ((operation_194_3706)>>(operation_194_2119));
            operation_194_3705 <= ((operation_194_3706)<<(operation_194_5557));
            operation_194_3707 <= ((operation_194_3708)&(operation_194_5557));
            operation_194_3708 <= ((operation_194_3710)>>(operation_194_2119));
            operation_194_3709 <= ((operation_194_3710)<<(operation_194_5557));
            operation_194_3713 <= ((operation_194_3784)^(operation_194_3813));
            operation_194_3716 <= ((operation_194_3782)^(operation_194_3811));
            operation_194_3719 <= ((operation_194_3780)^(operation_194_3809));
            operation_194_3722 <= ((operation_194_3778)^(operation_194_3807));
            operation_194_3724 <= ((operation_194_3740)^(operation_194_3813));
            operation_194_3726 <= ((operation_194_3738)^(operation_194_3809));
            operation_194_3728 <= ((operation_194_3735)^(operation_194_5577));
            operation_194_3730 <= ((operation_194_3185)^(operation_194_3734));
            operation_194_3732 <= ((operation_194_3184)^(operation_194_3733));
            operation_194_3738 <= ((operation_194_3739)^(operation_194_3780));
            operation_194_3739 <= ((operation_194_3779)^(operation_194_3810));
            operation_194_3740 <= ((operation_194_3741)^(operation_194_3784));
            operation_194_3741 <= ((operation_194_3783)^(operation_194_3814));
            operation_194_3743 <= ((operation_194_3814)^(operation_194_3784));
            operation_194_3745 <= ((operation_194_3813)^(operation_194_3783));
            operation_194_3747 <= ((operation_194_3812)^(operation_194_3782));
            operation_194_3749 <= ((operation_194_3811)^(operation_194_3781));
            operation_194_3751 <= ((operation_194_3810)^(operation_194_3780));
            operation_194_3753 <= ((operation_194_3809)^(operation_194_3779));
            operation_194_3755 <= ((operation_194_3808)^(operation_194_3778));
            operation_194_3757 <= ((operation_194_3807)^(operation_194_3777));
            operation_194_3759 <= ((operation_194_3775)^(operation_194_3811));
            operation_194_3761 <= ((operation_194_3773)^(operation_194_3807));
            operation_194_3763 <= ((operation_194_3246)^(operation_194_3770));
            operation_194_3773 <= ((operation_194_3774)^(operation_194_3778));
            operation_194_3774 <= ((operation_194_3777)^(operation_194_3808));
            operation_194_3775 <= ((operation_194_3776)^(operation_194_3782));
            operation_194_3776 <= ((operation_194_3781)^(operation_194_3812));
            operation_194_3788 <= ((operation_194_3305)^(operation_194_3803));
            operation_194_3790 <= ((operation_194_3304)^(operation_194_3801));
            operation_194_3805_latch <= (operation_194_3805);
            operation_194_3806_latch <= (operation_194_3806);
            operation_194_3815_latch <= (operation_194_3815);
            operation_194_3816_latch <= (operation_194_3816);
            operation_194_3817_latch <= (operation_194_3817);
            operation_194_3818_latch <= (operation_194_3818);
            operation_194_3819_latch <= (operation_194_3819);
            operation_194_3820_latch <= (operation_194_3820);
            operation_194_3821_latch <= (operation_194_3821);
            operation_194_3822_latch <= (operation_194_3822);
            operation_194_3823_latch <= (operation_194_3823);
            operation_194_3824_latch <= (operation_194_3824);
            operation_194_3825_latch <= (operation_194_3825);
            operation_194_3826_latch <= (operation_194_3826);
            operation_194_3827_latch <= (operation_194_3827);
            operation_194_3828_latch <= (operation_194_3828);
            operation_194_3829_latch <= (operation_194_3829);
            operation_194_3830_latch <= (operation_194_3830);
            operation_194_3831_latch <= (operation_194_3831);
            operation_194_3832_latch <= (operation_194_3832);
            operation_194_2987 <= ((operation_194_3008)^(operation_194_2988));
            operation_194_2991 <= ((operation_194_2559)^(operation_194_3015));
            operation_194_2993 <= ((operation_194_3014)^(operation_194_3147));
            operation_194_2995 <= ((operation_194_3013)^(operation_194_3246));
            operation_194_2997 <= ((operation_194_3012)^(operation_194_3087));
            operation_194_2999 <= ((operation_194_3011)^(operation_194_3146));
            operation_194_3001 <= ((operation_194_3010)^(operation_194_3015));
            operation_194_3003 <= ((operation_194_3009)^(operation_194_3086));
            operation_194_3005 <= ((operation_194_3007)^(operation_194_3006));
            operation_194_3017 <= ((operation_194_3354)^(operation_194_3065));
            operation_194_3019 <= ((operation_194_3355)^(operation_194_3064));
            operation_194_3021 <= ((operation_194_3352)^(operation_194_3063));
            operation_194_3023 <= ((operation_194_3353)^(operation_194_3062));
            operation_194_3025 <= ((operation_194_3350)^(operation_194_3061));
            operation_194_3027 <= ((operation_194_3351)^(operation_194_3060));
            operation_194_3029 <= ((operation_194_3348)^(operation_194_3059));
            operation_194_3031 <= ((operation_194_3349)^(operation_194_3058));
            operation_194_3033 <= ((operation_194_3057)^(operation_194_3305));
            operation_194_3035 <= ((operation_194_3056)^(operation_194_3304));
            operation_194_3037 <= ((operation_194_3055)^(operation_194_3185));
            operation_194_3039 <= ((operation_194_3054)^(operation_194_3184));
            operation_194_3041 <= ((operation_194_3053)^(operation_194_3117));
            operation_194_3043 <= ((operation_194_3052)^(operation_194_3116));
            operation_194_3045 <= ((operation_194_3051)^(operation_194_3050));
            operation_194_3047 <= ((operation_194_3049)^(operation_194_3048));
            operation_194_3067 <= ((operation_194_3385)^(operation_194_3095));
            operation_194_3069 <= ((operation_194_3384)^(operation_194_3094));
            operation_194_3071 <= ((operation_194_3383)^(operation_194_3093));
            operation_194_3073 <= ((operation_194_3382)^(operation_194_3092));
            operation_194_3075 <= ((operation_194_3381)^(operation_194_3091));
            operation_194_3077 <= ((operation_194_3380)^(operation_194_3090));
            operation_194_3079 <= ((operation_194_3379)^(operation_194_3089));
            operation_194_3081 <= ((operation_194_3378)^(operation_194_3088));
            operation_194_3083 <= ((operation_194_2586)^(operation_194_3087));
            operation_194_3085 <= ((operation_194_2577)^(operation_194_3086));
            operation_194_3097 <= ((operation_194_3125)^(operation_194_3249));
            operation_194_3099 <= ((operation_194_3124)^(operation_194_3249));
            operation_194_3101 <= ((operation_194_3123)^(operation_194_3308));
            operation_194_3103 <= ((operation_194_3122)^(operation_194_3308));
            operation_194_3105 <= ((operation_194_3121)^(operation_194_3248));
            operation_194_3107 <= ((operation_194_3120)^(operation_194_3248));
            operation_194_3109 <= ((operation_194_3119)^(operation_194_3307));
            operation_194_3111 <= ((operation_194_3118)^(operation_194_3307));
            operation_194_3113 <= ((operation_194_2621)^(operation_194_3117));
            operation_194_3115 <= ((operation_194_2619)^(operation_194_3116));
            operation_194_3127 <= ((operation_194_3155)^(operation_194_3249));
            operation_194_3129 <= ((operation_194_3154)^(operation_194_3249));
            operation_194_3131 <= ((operation_194_3153)^(operation_194_3308));
            operation_194_3133 <= ((operation_194_3152)^(operation_194_3308));
            operation_194_3135 <= ((operation_194_3151)^(operation_194_3248));
            operation_194_3137 <= ((operation_194_3150)^(operation_194_3248));
            operation_194_3139 <= ((operation_194_3149)^(operation_194_3307));
            operation_194_3141 <= ((operation_194_3148)^(operation_194_3307));
            operation_194_3143 <= ((operation_194_2658)^(operation_194_3147));
            operation_194_3145 <= ((operation_194_2657)^(operation_194_3146));
            operation_194_3157 <= ((operation_194_3216)^(operation_194_3158));
            operation_194_3158 <= ((operation_194_3214)*(operation_194_5597));
            operation_194_3160 <= ((operation_194_3212)^(operation_194_3161));
            operation_194_3161 <= ((operation_194_3210)*(operation_194_5597));
            operation_194_3163 <= ((operation_194_3208)^(operation_194_3164));
            operation_194_3164 <= ((operation_194_3206)*(operation_194_5597));
            operation_194_3166 <= ((operation_194_3204)^(operation_194_3167));
            operation_194_3167 <= ((operation_194_3202)*(operation_194_5597));
            operation_194_3169 <= ((operation_194_3200)^(operation_194_3170));
            operation_194_3170 <= ((operation_194_3198)*(operation_194_5597));
            operation_194_3172 <= ((operation_194_3196)^(operation_194_3173));
            operation_194_3173 <= ((operation_194_3194)*(operation_194_5597));
            operation_194_3175 <= ((operation_194_3192)^(operation_194_3176));
            operation_194_3176 <= ((operation_194_3190)*(operation_194_5597));
            operation_194_3178 <= ((operation_194_3188)^(operation_194_3179));
            operation_194_3179 <= ((operation_194_3186)*(operation_194_5597));
            operation_194_3181 <= ((operation_194_2688)^(operation_194_3185));
            operation_194_3183 <= ((operation_194_2687)^(operation_194_3184));
            operation_194_3186 <= ((operation_194_3187)&(operation_194_5557));
            operation_194_3187 <= ((operation_194_3189)>>(operation_194_2119));
            operation_194_3188 <= ((operation_194_3189)<<(operation_194_5557));
            operation_194_3190 <= ((operation_194_3191)&(operation_194_5557));
            operation_194_3191 <= ((operation_194_3193)>>(operation_194_2119));
            operation_194_3192 <= ((operation_194_3193)<<(operation_194_5557));
            operation_194_3194 <= ((operation_194_3195)&(operation_194_5557));
            operation_194_3195 <= ((operation_194_3197)>>(operation_194_2119));
            operation_194_3196 <= ((operation_194_3197)<<(operation_194_5557));
            operation_194_3198 <= ((operation_194_3199)&(operation_194_5557));
            operation_194_3199 <= ((operation_194_3201)>>(operation_194_2119));
            operation_194_3200 <= ((operation_194_3201)<<(operation_194_5557));
            operation_194_3202 <= ((operation_194_3203)&(operation_194_5557));
            operation_194_3203 <= ((operation_194_3205)>>(operation_194_2119));
            operation_194_3204 <= ((operation_194_3205)<<(operation_194_5557));
            operation_194_3206 <= ((operation_194_3207)&(operation_194_5557));
            operation_194_3207 <= ((operation_194_3209)>>(operation_194_2119));
            operation_194_3208 <= ((operation_194_3209)<<(operation_194_5557));
            operation_194_3210 <= ((operation_194_3211)&(operation_194_5557));
            operation_194_3211 <= ((operation_194_3213)>>(operation_194_2119));
            operation_194_3212 <= ((operation_194_3213)<<(operation_194_5557));
            operation_194_3214 <= ((operation_194_3215)&(operation_194_5557));
            operation_194_3215 <= ((operation_194_3217)>>(operation_194_2119));
            operation_194_3216 <= ((operation_194_3217)<<(operation_194_5557));
            operation_194_3219 <= ((operation_194_3280)^(operation_194_3220));
            operation_194_3220 <= ((operation_194_3278)*(operation_194_5597));
            operation_194_3222 <= ((operation_194_3276)^(operation_194_3223));
            operation_194_3223 <= ((operation_194_3274)*(operation_194_5597));
            operation_194_3225 <= ((operation_194_3272)^(operation_194_3226));
            operation_194_3226 <= ((operation_194_3270)*(operation_194_5597));
            operation_194_3228 <= ((operation_194_3268)^(operation_194_3229));
            operation_194_3229 <= ((operation_194_3266)*(operation_194_5597));
            operation_194_3231 <= ((operation_194_3264)^(operation_194_3232));
            operation_194_3232 <= ((operation_194_3262)*(operation_194_5597));
            operation_194_3234 <= ((operation_194_3260)^(operation_194_3235));
            operation_194_3235 <= ((operation_194_3258)*(operation_194_5597));
            operation_194_3237 <= ((operation_194_3256)^(operation_194_3238));
            operation_194_3238 <= ((operation_194_3254)*(operation_194_5597));
            operation_194_3240 <= ((operation_194_3252)^(operation_194_3241));
            operation_194_3241 <= ((operation_194_3250)*(operation_194_5597));
            operation_194_3243 <= ((operation_194_2718)^(operation_194_3247));
            operation_194_3245 <= ((operation_194_2717)^(operation_194_3246));
            operation_194_3250 <= ((operation_194_3251)&(operation_194_5557));
            operation_194_3251 <= ((operation_194_3253)>>(operation_194_2119));
            operation_194_3252 <= ((operation_194_3253)<<(operation_194_5557));
            operation_194_3254 <= ((operation_194_3255)&(operation_194_5557));
            operation_194_3255 <= ((operation_194_3257)>>(operation_194_2119));
            operation_194_3256 <= ((operation_194_3257)<<(operation_194_5557));
            operation_194_3258 <= ((operation_194_3259)&(operation_194_5557));
            operation_194_3259 <= ((operation_194_3261)>>(operation_194_2119));
            operation_194_3260 <= ((operation_194_3261)<<(operation_194_5557));
            operation_194_3262 <= ((operation_194_3263)&(operation_194_5557));
            operation_194_3263 <= ((operation_194_3265)>>(operation_194_2119));
            operation_194_3264 <= ((operation_194_3265)<<(operation_194_5557));
            operation_194_3266 <= ((operation_194_3267)&(operation_194_5557));
            operation_194_3267 <= ((operation_194_3269)>>(operation_194_2119));
            operation_194_3268 <= ((operation_194_3269)<<(operation_194_5557));
            operation_194_3270 <= ((operation_194_3271)&(operation_194_5557));
            operation_194_3271 <= ((operation_194_3273)>>(operation_194_2119));
            operation_194_3272 <= ((operation_194_3273)<<(operation_194_5557));
            operation_194_3274 <= ((operation_194_3275)&(operation_194_5557));
            operation_194_3275 <= ((operation_194_3277)>>(operation_194_2119));
            operation_194_3276 <= ((operation_194_3277)<<(operation_194_5557));
            operation_194_3278 <= ((operation_194_3279)&(operation_194_5557));
            operation_194_3279 <= ((operation_194_3281)>>(operation_194_2119));
            operation_194_3280 <= ((operation_194_3281)<<(operation_194_5557));
            operation_194_3284 <= ((operation_194_3355)^(operation_194_3384));
            operation_194_3287 <= ((operation_194_3353)^(operation_194_3382));
            operation_194_3290 <= ((operation_194_3351)^(operation_194_3380));
            operation_194_3293 <= ((operation_194_3349)^(operation_194_3378));
            operation_194_3295 <= ((operation_194_3311)^(operation_194_3384));
            operation_194_3297 <= ((operation_194_3309)^(operation_194_3380));
            operation_194_3299 <= ((operation_194_3306)^(operation_194_5572));
            operation_194_3301 <= ((operation_194_2756)^(operation_194_3305));
            operation_194_3303 <= ((operation_194_2755)^(operation_194_3304));
            operation_194_3309 <= ((operation_194_3310)^(operation_194_3351));
            operation_194_3310 <= ((operation_194_3350)^(operation_194_3381));
            operation_194_3311 <= ((operation_194_3312)^(operation_194_3355));
            operation_194_3312 <= ((operation_194_3354)^(operation_194_3385));
            operation_194_3314 <= ((operation_194_3385)^(operation_194_3355));
            operation_194_3316 <= ((operation_194_3384)^(operation_194_3354));
            operation_194_3318 <= ((operation_194_3383)^(operation_194_3353));
            operation_194_3320 <= ((operation_194_3382)^(operation_194_3352));
            operation_194_3322 <= ((operation_194_3381)^(operation_194_3351));
            operation_194_3324 <= ((operation_194_3380)^(operation_194_3350));
            operation_194_3326 <= ((operation_194_3379)^(operation_194_3349));
            operation_194_3328 <= ((operation_194_3378)^(operation_194_3348));
            operation_194_3330 <= ((operation_194_3346)^(operation_194_3382));
            operation_194_3332 <= ((operation_194_3344)^(operation_194_3378));
            operation_194_3334 <= ((operation_194_2817)^(operation_194_3341));
            operation_194_3344 <= ((operation_194_3345)^(operation_194_3349));
            operation_194_3345 <= ((operation_194_3348)^(operation_194_3379));
            operation_194_3346 <= ((operation_194_3347)^(operation_194_3353));
            operation_194_3347 <= ((operation_194_3352)^(operation_194_3383));
            operation_194_3359 <= ((operation_194_2876)^(operation_194_3374));
            operation_194_3361 <= ((operation_194_2875)^(operation_194_3372));
            operation_194_3376_latch <= (operation_194_3376);
            operation_194_3377_latch <= (operation_194_3377);
            operation_194_3386_latch <= (operation_194_3386);
            operation_194_3387_latch <= (operation_194_3387);
            operation_194_3388_latch <= (operation_194_3388);
            operation_194_3389_latch <= (operation_194_3389);
            operation_194_3390_latch <= (operation_194_3390);
            operation_194_3391_latch <= (operation_194_3391);
            operation_194_3392_latch <= (operation_194_3392);
            operation_194_3393_latch <= (operation_194_3393);
            operation_194_3394_latch <= (operation_194_3394);
            operation_194_3395_latch <= (operation_194_3395);
            operation_194_3396_latch <= (operation_194_3396);
            operation_194_3397_latch <= (operation_194_3397);
            operation_194_3398_latch <= (operation_194_3398);
            operation_194_3399_latch <= (operation_194_3399);
            operation_194_3400_latch <= (operation_194_3400);
            operation_194_3401_latch <= (operation_194_3401);
            operation_194_3402_latch <= (operation_194_3402);
            operation_194_3403_latch <= (operation_194_3403);
            operation_194_2558 <= ((operation_194_2579)^(operation_194_2559));
            operation_194_2562 <= ((operation_194_2130)^(operation_194_2586));
            operation_194_2564 <= ((operation_194_2585)^(operation_194_2718));
            operation_194_2566 <= ((operation_194_2584)^(operation_194_2817));
            operation_194_2568 <= ((operation_194_2583)^(operation_194_2658));
            operation_194_2570 <= ((operation_194_2582)^(operation_194_2717));
            operation_194_2572 <= ((operation_194_2581)^(operation_194_2586));
            operation_194_2574 <= ((operation_194_2580)^(operation_194_2657));
            operation_194_2576 <= ((operation_194_2578)^(operation_194_2577));
            operation_194_2588 <= ((operation_194_2925)^(operation_194_2636));
            operation_194_2590 <= ((operation_194_2926)^(operation_194_2635));
            operation_194_2592 <= ((operation_194_2923)^(operation_194_2634));
            operation_194_2594 <= ((operation_194_2924)^(operation_194_2633));
            operation_194_2596 <= ((operation_194_2921)^(operation_194_2632));
            operation_194_2598 <= ((operation_194_2922)^(operation_194_2631));
            operation_194_2600 <= ((operation_194_2919)^(operation_194_2630));
            operation_194_2602 <= ((operation_194_2920)^(operation_194_2629));
            operation_194_2604 <= ((operation_194_2628)^(operation_194_2876));
            operation_194_2606 <= ((operation_194_2627)^(operation_194_2875));
            operation_194_2608 <= ((operation_194_2626)^(operation_194_2756));
            operation_194_2610 <= ((operation_194_2625)^(operation_194_2755));
            operation_194_2612 <= ((operation_194_2624)^(operation_194_2688));
            operation_194_2614 <= ((operation_194_2623)^(operation_194_2687));
            operation_194_2616 <= ((operation_194_2622)^(operation_194_2621));
            operation_194_2618 <= ((operation_194_2620)^(operation_194_2619));
            operation_194_2638 <= ((operation_194_2956)^(operation_194_2666));
            operation_194_2640 <= ((operation_194_2955)^(operation_194_2665));
            operation_194_2642 <= ((operation_194_2954)^(operation_194_2664));
            operation_194_2644 <= ((operation_194_2953)^(operation_194_2663));
            operation_194_2646 <= ((operation_194_2952)^(operation_194_2662));
            operation_194_2648 <= ((operation_194_2951)^(operation_194_2661));
            operation_194_2650 <= ((operation_194_2950)^(operation_194_2660));
            operation_194_2652 <= ((operation_194_2949)^(operation_194_2659));
            operation_194_2654 <= ((operation_194_2157)^(operation_194_2658));
            operation_194_2656 <= ((operation_194_2148)^(operation_194_2657));
            operation_194_2668 <= ((operation_194_2696)^(operation_194_2820));
            operation_194_2670 <= ((operation_194_2695)^(operation_194_2820));
            operation_194_2672 <= ((operation_194_2694)^(operation_194_2879));
            operation_194_2674 <= ((operation_194_2693)^(operation_194_2879));
            operation_194_2676 <= ((operation_194_2692)^(operation_194_2819));
            operation_194_2678 <= ((operation_194_2691)^(operation_194_2819));
            operation_194_2680 <= ((operation_194_2690)^(operation_194_2878));
            operation_194_2682 <= ((operation_194_2689)^(operation_194_2878));
            operation_194_2684 <= ((operation_194_2192)^(operation_194_2688));
            operation_194_2686 <= ((operation_194_2190)^(operation_194_2687));
            operation_194_2698 <= ((operation_194_2726)^(operation_194_2820));
            operation_194_2700 <= ((operation_194_2725)^(operation_194_2820));
            operation_194_2702 <= ((operation_194_2724)^(operation_194_2879));
            operation_194_2704 <= ((operation_194_2723)^(operation_194_2879));
            operation_194_2706 <= ((operation_194_2722)^(operation_194_2819));
            operation_194_2708 <= ((operation_194_2721)^(operation_194_2819));
            operation_194_2710 <= ((operation_194_2720)^(operation_194_2878));
            operation_194_2712 <= ((operation_194_2719)^(operation_194_2878));
            operation_194_2714 <= ((operation_194_2229)^(operation_194_2718));
            operation_194_2716 <= ((operation_194_2228)^(operation_194_2717));
            operation_194_2728 <= ((operation_194_2787)^(operation_194_2729));
            operation_194_2729 <= ((operation_194_2785)*(operation_194_5597));
            operation_194_2731 <= ((operation_194_2783)^(operation_194_2732));
            operation_194_2732 <= ((operation_194_2781)*(operation_194_5597));
            operation_194_2734 <= ((operation_194_2779)^(operation_194_2735));
            operation_194_2735 <= ((operation_194_2777)*(operation_194_5597));
            operation_194_2737 <= ((operation_194_2775)^(operation_194_2738));
            operation_194_2738 <= ((operation_194_2773)*(operation_194_5597));
            operation_194_2740 <= ((operation_194_2771)^(operation_194_2741));
            operation_194_2741 <= ((operation_194_2769)*(operation_194_5597));
            operation_194_2743 <= ((operation_194_2767)^(operation_194_2744));
            operation_194_2744 <= ((operation_194_2765)*(operation_194_5597));
            operation_194_2746 <= ((operation_194_2763)^(operation_194_2747));
            operation_194_2747 <= ((operation_194_2761)*(operation_194_5597));
            operation_194_2749 <= ((operation_194_2759)^(operation_194_2750));
            operation_194_2750 <= ((operation_194_2757)*(operation_194_5597));
            operation_194_2752 <= ((operation_194_2259)^(operation_194_2756));
            operation_194_2754 <= ((operation_194_2258)^(operation_194_2755));
            operation_194_2757 <= ((operation_194_2758)&(operation_194_5557));
            operation_194_2758 <= ((operation_194_2760)>>(operation_194_2119));
            operation_194_2759 <= ((operation_194_2760)<<(operation_194_5557));
            operation_194_2761 <= ((operation_194_2762)&(operation_194_5557));
            operation_194_2762 <= ((operation_194_2764)>>(operation_194_2119));
            operation_194_2763 <= ((operation_194_2764)<<(operation_194_5557));
            operation_194_2765 <= ((operation_194_2766)&(operation_194_5557));
            operation_194_2766 <= ((operation_194_2768)>>(operation_194_2119));
            operation_194_2767 <= ((operation_194_2768)<<(operation_194_5557));
            operation_194_2769 <= ((operation_194_2770)&(operation_194_5557));
            operation_194_2770 <= ((operation_194_2772)>>(operation_194_2119));
            operation_194_2771 <= ((operation_194_2772)<<(operation_194_5557));
            operation_194_2773 <= ((operation_194_2774)&(operation_194_5557));
            operation_194_2774 <= ((operation_194_2776)>>(operation_194_2119));
            operation_194_2775 <= ((operation_194_2776)<<(operation_194_5557));
            operation_194_2777 <= ((operation_194_2778)&(operation_194_5557));
            operation_194_2778 <= ((operation_194_2780)>>(operation_194_2119));
            operation_194_2779 <= ((operation_194_2780)<<(operation_194_5557));
            operation_194_2781 <= ((operation_194_2782)&(operation_194_5557));
            operation_194_2782 <= ((operation_194_2784)>>(operation_194_2119));
            operation_194_2783 <= ((operation_194_2784)<<(operation_194_5557));
            operation_194_2785 <= ((operation_194_2786)&(operation_194_5557));
            operation_194_2786 <= ((operation_194_2788)>>(operation_194_2119));
            operation_194_2787 <= ((operation_194_2788)<<(operation_194_5557));
            operation_194_2790 <= ((operation_194_2851)^(operation_194_2791));
            operation_194_2791 <= ((operation_194_2849)*(operation_194_5597));
            operation_194_2793 <= ((operation_194_2847)^(operation_194_2794));
            operation_194_2794 <= ((operation_194_2845)*(operation_194_5597));
            operation_194_2796 <= ((operation_194_2843)^(operation_194_2797));
            operation_194_2797 <= ((operation_194_2841)*(operation_194_5597));
            operation_194_2799 <= ((operation_194_2839)^(operation_194_2800));
            operation_194_2800 <= ((operation_194_2837)*(operation_194_5597));
            operation_194_2802 <= ((operation_194_2835)^(operation_194_2803));
            operation_194_2803 <= ((operation_194_2833)*(operation_194_5597));
            operation_194_2805 <= ((operation_194_2831)^(operation_194_2806));
            operation_194_2806 <= ((operation_194_2829)*(operation_194_5597));
            operation_194_2808 <= ((operation_194_2827)^(operation_194_2809));
            operation_194_2809 <= ((operation_194_2825)*(operation_194_5597));
            operation_194_2811 <= ((operation_194_2823)^(operation_194_2812));
            operation_194_2812 <= ((operation_194_2821)*(operation_194_5597));
            operation_194_2814 <= ((operation_194_2289)^(operation_194_2818));
            operation_194_2816 <= ((operation_194_2288)^(operation_194_2817));
            operation_194_2821 <= ((operation_194_2822)&(operation_194_5557));
            operation_194_2822 <= ((operation_194_2824)>>(operation_194_2119));
            operation_194_2823 <= ((operation_194_2824)<<(operation_194_5557));
            operation_194_2825 <= ((operation_194_2826)&(operation_194_5557));
            operation_194_2826 <= ((operation_194_2828)>>(operation_194_2119));
            operation_194_2827 <= ((operation_194_2828)<<(operation_194_5557));
            operation_194_2829 <= ((operation_194_2830)&(operation_194_5557));
            operation_194_2830 <= ((operation_194_2832)>>(operation_194_2119));
            operation_194_2831 <= ((operation_194_2832)<<(operation_194_5557));
            operation_194_2833 <= ((operation_194_2834)&(operation_194_5557));
            operation_194_2834 <= ((operation_194_2836)>>(operation_194_2119));
            operation_194_2835 <= ((operation_194_2836)<<(operation_194_5557));
            operation_194_2837 <= ((operation_194_2838)&(operation_194_5557));
            operation_194_2838 <= ((operation_194_2840)>>(operation_194_2119));
            operation_194_2839 <= ((operation_194_2840)<<(operation_194_5557));
            operation_194_2841 <= ((operation_194_2842)&(operation_194_5557));
            operation_194_2842 <= ((operation_194_2844)>>(operation_194_2119));
            operation_194_2843 <= ((operation_194_2844)<<(operation_194_5557));
            operation_194_2845 <= ((operation_194_2846)&(operation_194_5557));
            operation_194_2846 <= ((operation_194_2848)>>(operation_194_2119));
            operation_194_2847 <= ((operation_194_2848)<<(operation_194_5557));
            operation_194_2849 <= ((operation_194_2850)&(operation_194_5557));
            operation_194_2850 <= ((operation_194_2852)>>(operation_194_2119));
            operation_194_2851 <= ((operation_194_2852)<<(operation_194_5557));
            operation_194_2855 <= ((operation_194_2926)^(operation_194_2955));
            operation_194_2858 <= ((operation_194_2924)^(operation_194_2953));
            operation_194_2861 <= ((operation_194_2922)^(operation_194_2951));
            operation_194_2864 <= ((operation_194_2920)^(operation_194_2949));
            operation_194_2866 <= ((operation_194_2882)^(operation_194_2955));
            operation_194_2868 <= ((operation_194_2880)^(operation_194_2951));
            operation_194_2870 <= ((operation_194_2877)^(operation_194_5567));
            operation_194_2872 <= ((operation_194_2327)^(operation_194_2876));
            operation_194_2874 <= ((operation_194_2326)^(operation_194_2875));
            operation_194_2880 <= ((operation_194_2881)^(operation_194_2922));
            operation_194_2881 <= ((operation_194_2921)^(operation_194_2952));
            operation_194_2882 <= ((operation_194_2883)^(operation_194_2926));
            operation_194_2883 <= ((operation_194_2925)^(operation_194_2956));
            operation_194_2885 <= ((operation_194_2956)^(operation_194_2926));
            operation_194_2887 <= ((operation_194_2955)^(operation_194_2925));
            operation_194_2889 <= ((operation_194_2954)^(operation_194_2924));
            operation_194_2891 <= ((operation_194_2953)^(operation_194_2923));
            operation_194_2893 <= ((operation_194_2952)^(operation_194_2922));
            operation_194_2895 <= ((operation_194_2951)^(operation_194_2921));
            operation_194_2897 <= ((operation_194_2950)^(operation_194_2920));
            operation_194_2899 <= ((operation_194_2949)^(operation_194_2919));
            operation_194_2901 <= ((operation_194_2917)^(operation_194_2953));
            operation_194_2903 <= ((operation_194_2915)^(operation_194_2949));
            operation_194_2905 <= ((operation_194_2388)^(operation_194_2912));
            operation_194_2915 <= ((operation_194_2916)^(operation_194_2920));
            operation_194_2916 <= ((operation_194_2919)^(operation_194_2950));
            operation_194_2917 <= ((operation_194_2918)^(operation_194_2924));
            operation_194_2918 <= ((operation_194_2923)^(operation_194_2954));
            operation_194_2930 <= ((operation_194_2447)^(operation_194_2945));
            operation_194_2932 <= ((operation_194_2446)^(operation_194_2943));
            operation_194_2947_latch <= (operation_194_2947);
            operation_194_2948_latch <= (operation_194_2948);
            operation_194_2957_latch <= (operation_194_2957);
            operation_194_2958_latch <= (operation_194_2958);
            operation_194_2959_latch <= (operation_194_2959);
            operation_194_2960_latch <= (operation_194_2960);
            operation_194_2961_latch <= (operation_194_2961);
            operation_194_2962_latch <= (operation_194_2962);
            operation_194_2963_latch <= (operation_194_2963);
            operation_194_2964_latch <= (operation_194_2964);
            operation_194_2965_latch <= (operation_194_2965);
            operation_194_2966_latch <= (operation_194_2966);
            operation_194_2967_latch <= (operation_194_2967);
            operation_194_2968_latch <= (operation_194_2968);
            operation_194_2969_latch <= (operation_194_2969);
            operation_194_2970_latch <= (operation_194_2970);
            operation_194_2971_latch <= (operation_194_2971);
            operation_194_2972_latch <= (operation_194_2972);
            operation_194_2973_latch <= (operation_194_2973);
            operation_194_2974_latch <= (operation_194_2974);
            operation_194_2129 <= ((operation_194_2150)^(operation_194_2130));
            operation_194_2133 <= ((operation_194_1701)^(operation_194_2157));
            operation_194_2135 <= ((operation_194_2156)^(operation_194_2289));
            operation_194_2137 <= ((operation_194_2155)^(operation_194_2388));
            operation_194_2139 <= ((operation_194_2154)^(operation_194_2229));
            operation_194_2141 <= ((operation_194_2153)^(operation_194_2288));
            operation_194_2143 <= ((operation_194_2152)^(operation_194_2157));
            operation_194_2145 <= ((operation_194_2151)^(operation_194_2228));
            operation_194_2147 <= ((operation_194_2149)^(operation_194_2148));
            operation_194_2159 <= ((operation_194_2496)^(operation_194_2207));
            operation_194_2161 <= ((operation_194_2497)^(operation_194_2206));
            operation_194_2163 <= ((operation_194_2494)^(operation_194_2205));
            operation_194_2165 <= ((operation_194_2495)^(operation_194_2204));
            operation_194_2167 <= ((operation_194_2492)^(operation_194_2203));
            operation_194_2169 <= ((operation_194_2493)^(operation_194_2202));
            operation_194_2171 <= ((operation_194_2490)^(operation_194_2201));
            operation_194_2173 <= ((operation_194_2491)^(operation_194_2200));
            operation_194_2175 <= ((operation_194_2199)^(operation_194_2447));
            operation_194_2177 <= ((operation_194_2198)^(operation_194_2446));
            operation_194_2179 <= ((operation_194_2197)^(operation_194_2327));
            operation_194_2181 <= ((operation_194_2196)^(operation_194_2326));
            operation_194_2183 <= ((operation_194_2195)^(operation_194_2259));
            operation_194_2185 <= ((operation_194_2194)^(operation_194_2258));
            operation_194_2187 <= ((operation_194_2193)^(operation_194_2192));
            operation_194_2189 <= ((operation_194_2191)^(operation_194_2190));
            operation_194_2209 <= ((operation_194_2527)^(operation_194_2237));
            operation_194_2211 <= ((operation_194_2526)^(operation_194_2236));
            operation_194_2213 <= ((operation_194_2525)^(operation_194_2235));
            operation_194_2215 <= ((operation_194_2524)^(operation_194_2234));
            operation_194_2217 <= ((operation_194_2523)^(operation_194_2233));
            operation_194_2219 <= ((operation_194_2522)^(operation_194_2232));
            operation_194_2221 <= ((operation_194_2521)^(operation_194_2231));
            operation_194_2223 <= ((operation_194_2520)^(operation_194_2230));
            operation_194_2225 <= ((operation_194_1728)^(operation_194_2229));
            operation_194_2227 <= ((operation_194_1719)^(operation_194_2228));
            operation_194_2239 <= ((operation_194_2267)^(operation_194_2391));
            operation_194_2241 <= ((operation_194_2266)^(operation_194_2391));
            operation_194_2243 <= ((operation_194_2265)^(operation_194_2450));
            operation_194_2245 <= ((operation_194_2264)^(operation_194_2450));
            operation_194_2247 <= ((operation_194_2263)^(operation_194_2390));
            operation_194_2249 <= ((operation_194_2262)^(operation_194_2390));
            operation_194_2251 <= ((operation_194_2261)^(operation_194_2449));
            operation_194_2253 <= ((operation_194_2260)^(operation_194_2449));
            operation_194_2255 <= ((operation_194_1763)^(operation_194_2259));
            operation_194_2257 <= ((operation_194_1761)^(operation_194_2258));
            operation_194_2269 <= ((operation_194_2297)^(operation_194_2391));
            operation_194_2271 <= ((operation_194_2296)^(operation_194_2391));
            operation_194_2273 <= ((operation_194_2295)^(operation_194_2450));
            operation_194_2275 <= ((operation_194_2294)^(operation_194_2450));
            operation_194_2277 <= ((operation_194_2293)^(operation_194_2390));
            operation_194_2279 <= ((operation_194_2292)^(operation_194_2390));
            operation_194_2281 <= ((operation_194_2291)^(operation_194_2449));
            operation_194_2283 <= ((operation_194_2290)^(operation_194_2449));
            operation_194_2285 <= ((operation_194_1800)^(operation_194_2289));
            operation_194_2287 <= ((operation_194_1799)^(operation_194_2288));
            operation_194_2299 <= ((operation_194_2358)^(operation_194_2300));
            operation_194_2300 <= ((operation_194_2356)*(operation_194_5597));
            operation_194_2302 <= ((operation_194_2354)^(operation_194_2303));
            operation_194_2303 <= ((operation_194_2352)*(operation_194_5597));
            operation_194_2305 <= ((operation_194_2350)^(operation_194_2306));
            operation_194_2306 <= ((operation_194_2348)*(operation_194_5597));
            operation_194_2308 <= ((operation_194_2346)^(operation_194_2309));
            operation_194_2309 <= ((operation_194_2344)*(operation_194_5597));
            operation_194_2311 <= ((operation_194_2342)^(operation_194_2312));
            operation_194_2312 <= ((operation_194_2340)*(operation_194_5597));
            operation_194_2314 <= ((operation_194_2338)^(operation_194_2315));
            operation_194_2315 <= ((operation_194_2336)*(operation_194_5597));
            operation_194_2317 <= ((operation_194_2334)^(operation_194_2318));
            operation_194_2318 <= ((operation_194_2332)*(operation_194_5597));
            operation_194_2320 <= ((operation_194_2330)^(operation_194_2321));
            operation_194_2321 <= ((operation_194_2328)*(operation_194_5597));
            operation_194_2323 <= ((operation_194_1830)^(operation_194_2327));
            operation_194_2325 <= ((operation_194_1829)^(operation_194_2326));
            operation_194_2328 <= ((operation_194_2329)&(operation_194_5557));
            operation_194_2329 <= ((operation_194_2331)>>(operation_194_2119));
            operation_194_2330 <= ((operation_194_2331)<<(operation_194_5557));
            operation_194_2332 <= ((operation_194_2333)&(operation_194_5557));
            operation_194_2333 <= ((operation_194_2335)>>(operation_194_2119));
            operation_194_2334 <= ((operation_194_2335)<<(operation_194_5557));
            operation_194_2336 <= ((operation_194_2337)&(operation_194_5557));
            operation_194_2337 <= ((operation_194_2339)>>(operation_194_2119));
            operation_194_2338 <= ((operation_194_2339)<<(operation_194_5557));
            operation_194_2340 <= ((operation_194_2341)&(operation_194_5557));
            operation_194_2341 <= ((operation_194_2343)>>(operation_194_2119));
            operation_194_2342 <= ((operation_194_2343)<<(operation_194_5557));
            operation_194_2344 <= ((operation_194_2345)&(operation_194_5557));
            operation_194_2345 <= ((operation_194_2347)>>(operation_194_2119));
            operation_194_2346 <= ((operation_194_2347)<<(operation_194_5557));
            operation_194_2348 <= ((operation_194_2349)&(operation_194_5557));
            operation_194_2349 <= ((operation_194_2351)>>(operation_194_2119));
            operation_194_2350 <= ((operation_194_2351)<<(operation_194_5557));
            operation_194_2352 <= ((operation_194_2353)&(operation_194_5557));
            operation_194_2353 <= ((operation_194_2355)>>(operation_194_2119));
            operation_194_2354 <= ((operation_194_2355)<<(operation_194_5557));
            operation_194_2356 <= ((operation_194_2357)&(operation_194_5557));
            operation_194_2357 <= ((operation_194_2359)>>(operation_194_2119));
            operation_194_2358 <= ((operation_194_2359)<<(operation_194_5557));
            operation_194_2361 <= ((operation_194_2422)^(operation_194_2362));
            operation_194_2362 <= ((operation_194_2420)*(operation_194_5597));
            operation_194_2364 <= ((operation_194_2418)^(operation_194_2365));
            operation_194_2365 <= ((operation_194_2416)*(operation_194_5597));
            operation_194_2367 <= ((operation_194_2414)^(operation_194_2368));
            operation_194_2368 <= ((operation_194_2412)*(operation_194_5597));
            operation_194_2370 <= ((operation_194_2410)^(operation_194_2371));
            operation_194_2371 <= ((operation_194_2408)*(operation_194_5597));
            operation_194_2373 <= ((operation_194_2406)^(operation_194_2374));
            operation_194_2374 <= ((operation_194_2404)*(operation_194_5597));
            operation_194_2376 <= ((operation_194_2402)^(operation_194_2377));
            operation_194_2377 <= ((operation_194_2400)*(operation_194_5597));
            operation_194_2379 <= ((operation_194_2398)^(operation_194_2380));
            operation_194_2380 <= ((operation_194_2396)*(operation_194_5597));
            operation_194_2382 <= ((operation_194_2394)^(operation_194_2383));
            operation_194_2383 <= ((operation_194_2392)*(operation_194_5597));
            operation_194_2385 <= ((operation_194_1860)^(operation_194_2389));
            operation_194_2387 <= ((operation_194_1859)^(operation_194_2388));
            operation_194_2392 <= ((operation_194_2393)&(operation_194_5557));
            operation_194_2393 <= ((operation_194_2395)>>(operation_194_2119));
            operation_194_2394 <= ((operation_194_2395)<<(operation_194_5557));
            operation_194_2396 <= ((operation_194_2397)&(operation_194_5557));
            operation_194_2397 <= ((operation_194_2399)>>(operation_194_2119));
            operation_194_2398 <= ((operation_194_2399)<<(operation_194_5557));
            operation_194_2400 <= ((operation_194_2401)&(operation_194_5557));
            operation_194_2401 <= ((operation_194_2403)>>(operation_194_2119));
            operation_194_2402 <= ((operation_194_2403)<<(operation_194_5557));
            operation_194_2404 <= ((operation_194_2405)&(operation_194_5557));
            operation_194_2405 <= ((operation_194_2407)>>(operation_194_2119));
            operation_194_2406 <= ((operation_194_2407)<<(operation_194_5557));
            operation_194_2408 <= ((operation_194_2409)&(operation_194_5557));
            operation_194_2409 <= ((operation_194_2411)>>(operation_194_2119));
            operation_194_2410 <= ((operation_194_2411)<<(operation_194_5557));
            operation_194_2412 <= ((operation_194_2413)&(operation_194_5557));
            operation_194_2413 <= ((operation_194_2415)>>(operation_194_2119));
            operation_194_2414 <= ((operation_194_2415)<<(operation_194_5557));
            operation_194_2416 <= ((operation_194_2417)&(operation_194_5557));
            operation_194_2417 <= ((operation_194_2419)>>(operation_194_2119));
            operation_194_2418 <= ((operation_194_2419)<<(operation_194_5557));
            operation_194_2420 <= ((operation_194_2421)&(operation_194_5557));
            operation_194_2421 <= ((operation_194_2423)>>(operation_194_2119));
            operation_194_2422 <= ((operation_194_2423)<<(operation_194_5557));
            operation_194_2426 <= ((operation_194_2497)^(operation_194_2526));
            operation_194_2429 <= ((operation_194_2495)^(operation_194_2524));
            operation_194_2432 <= ((operation_194_2493)^(operation_194_2522));
            operation_194_2435 <= ((operation_194_2491)^(operation_194_2520));
            operation_194_2437 <= ((operation_194_2453)^(operation_194_2526));
            operation_194_2439 <= ((operation_194_2451)^(operation_194_2522));
            operation_194_2441 <= ((operation_194_2448)^(operation_194_5562));
            operation_194_2443 <= ((operation_194_1898)^(operation_194_2447));
            operation_194_2445 <= ((operation_194_1897)^(operation_194_2446));
            operation_194_2451 <= ((operation_194_2452)^(operation_194_2493));
            operation_194_2452 <= ((operation_194_2492)^(operation_194_2523));
            operation_194_2453 <= ((operation_194_2454)^(operation_194_2497));
            operation_194_2454 <= ((operation_194_2496)^(operation_194_2527));
            operation_194_2456 <= ((operation_194_2527)^(operation_194_2497));
            operation_194_2458 <= ((operation_194_2526)^(operation_194_2496));
            operation_194_2460 <= ((operation_194_2525)^(operation_194_2495));
            operation_194_2462 <= ((operation_194_2524)^(operation_194_2494));
            operation_194_2464 <= ((operation_194_2523)^(operation_194_2493));
            operation_194_2466 <= ((operation_194_2522)^(operation_194_2492));
            operation_194_2468 <= ((operation_194_2521)^(operation_194_2491));
            operation_194_2470 <= ((operation_194_2520)^(operation_194_2490));
            operation_194_2472 <= ((operation_194_2488)^(operation_194_2524));
            operation_194_2474 <= ((operation_194_2486)^(operation_194_2520));
            operation_194_2476 <= ((operation_194_1959)^(operation_194_2483));
            operation_194_2486 <= ((operation_194_2487)^(operation_194_2491));
            operation_194_2487 <= ((operation_194_2490)^(operation_194_2521));
            operation_194_2488 <= ((operation_194_2489)^(operation_194_2495));
            operation_194_2489 <= ((operation_194_2494)^(operation_194_2525));
            operation_194_2501 <= ((operation_194_2018)^(operation_194_2516));
            operation_194_2503 <= ((operation_194_2017)^(operation_194_2514));
            operation_194_2518_latch <= (operation_194_2518);
            operation_194_2519_latch <= (operation_194_2519);
            operation_194_2528_latch <= (operation_194_2528);
            operation_194_2529_latch <= (operation_194_2529);
            operation_194_2530_latch <= (operation_194_2530);
            operation_194_2531_latch <= (operation_194_2531);
            operation_194_2532_latch <= (operation_194_2532);
            operation_194_2533_latch <= (operation_194_2533);
            operation_194_2534_latch <= (operation_194_2534);
            operation_194_2535_latch <= (operation_194_2535);
            operation_194_2536_latch <= (operation_194_2536);
            operation_194_2537_latch <= (operation_194_2537);
            operation_194_2538_latch <= (operation_194_2538);
            operation_194_2539_latch <= (operation_194_2539);
            operation_194_2540_latch <= (operation_194_2540);
            operation_194_2541_latch <= (operation_194_2541);
            operation_194_2542_latch <= (operation_194_2542);
            operation_194_2543_latch <= (operation_194_2543);
            operation_194_2544_latch <= (operation_194_2544);
            operation_194_2545_latch <= (operation_194_2545);
            operation_194_1700 <= ((operation_194_1721)^(operation_194_1701));
            operation_194_1704 <= ((operation_194_101)^(operation_194_1728));
            operation_194_1706 <= ((operation_194_1727)^(operation_194_1860));
            operation_194_1708 <= ((operation_194_1726)^(operation_194_1959));
            operation_194_1710 <= ((operation_194_1725)^(operation_194_1800));
            operation_194_1712 <= ((operation_194_1724)^(operation_194_1859));
            operation_194_1714 <= ((operation_194_1723)^(operation_194_1728));
            operation_194_1716 <= ((operation_194_1722)^(operation_194_1799));
            operation_194_1718 <= ((operation_194_1720)^(operation_194_1719));
            operation_194_1730 <= ((operation_194_2067)^(operation_194_1778));
            operation_194_1732 <= ((operation_194_2068)^(operation_194_1777));
            operation_194_1734 <= ((operation_194_2065)^(operation_194_1776));
            operation_194_1736 <= ((operation_194_2066)^(operation_194_1775));
            operation_194_1738 <= ((operation_194_2063)^(operation_194_1774));
            operation_194_1740 <= ((operation_194_2064)^(operation_194_1773));
            operation_194_1742 <= ((operation_194_2061)^(operation_194_1772));
            operation_194_1744 <= ((operation_194_2062)^(operation_194_1771));
            operation_194_1746 <= ((operation_194_1770)^(operation_194_2018));
            operation_194_1748 <= ((operation_194_1769)^(operation_194_2017));
            operation_194_1750 <= ((operation_194_1768)^(operation_194_1898));
            operation_194_1752 <= ((operation_194_1767)^(operation_194_1897));
            operation_194_1754 <= ((operation_194_1766)^(operation_194_1830));
            operation_194_1756 <= ((operation_194_1765)^(operation_194_1829));
            operation_194_1758 <= ((operation_194_1764)^(operation_194_1763));
            operation_194_1760 <= ((operation_194_1762)^(operation_194_1761));
            operation_194_1780 <= ((operation_194_2098)^(operation_194_1808));
            operation_194_1782 <= ((operation_194_2097)^(operation_194_1807));
            operation_194_1784 <= ((operation_194_2096)^(operation_194_1806));
            operation_194_1786 <= ((operation_194_2095)^(operation_194_1805));
            operation_194_1788 <= ((operation_194_2094)^(operation_194_1804));
            operation_194_1790 <= ((operation_194_2093)^(operation_194_1803));
            operation_194_1792 <= ((operation_194_2092)^(operation_194_1802));
            operation_194_1794 <= ((operation_194_2091)^(operation_194_1801));
            operation_194_1796 <= ((operation_194_69)^(operation_194_1800));
            operation_194_1798 <= ((operation_194_117)^(operation_194_1799));
            operation_194_1810 <= ((operation_194_1838)^(operation_194_1962));
            operation_194_1812 <= ((operation_194_1837)^(operation_194_1962));
            operation_194_1814 <= ((operation_194_1836)^(operation_194_2021));
            operation_194_1816 <= ((operation_194_1835)^(operation_194_2021));
            operation_194_1818 <= ((operation_194_1834)^(operation_194_1961));
            operation_194_1820 <= ((operation_194_1833)^(operation_194_1961));
            operation_194_1822 <= ((operation_194_1832)^(operation_194_2020));
            operation_194_1824 <= ((operation_194_1831)^(operation_194_2020));
            operation_194_1826 <= ((operation_194_109)^(operation_194_1830));
            operation_194_1828 <= ((operation_194_125)^(operation_194_1829));
            operation_194_1840 <= ((operation_194_1868)^(operation_194_1962));
            operation_194_1842 <= ((operation_194_1867)^(operation_194_1962));
            operation_194_1844 <= ((operation_194_1866)^(operation_194_2021));
            operation_194_1846 <= ((operation_194_1865)^(operation_194_2021));
            operation_194_1848 <= ((operation_194_1864)^(operation_194_1961));
            operation_194_1850 <= ((operation_194_1863)^(operation_194_1961));
            operation_194_1852 <= ((operation_194_1862)^(operation_194_2020));
            operation_194_1854 <= ((operation_194_1861)^(operation_194_2020));
            operation_194_1856 <= ((operation_194_37)^(operation_194_1860));
            operation_194_1858 <= ((operation_194_85)^(operation_194_1859));
            operation_194_1870 <= ((operation_194_1929)^(operation_194_1871));
            operation_194_1871 <= ((operation_194_1927)*(operation_194_5597));
            operation_194_1873 <= ((operation_194_1925)^(operation_194_1874));
            operation_194_1874 <= ((operation_194_1923)*(operation_194_5597));
            operation_194_1876 <= ((operation_194_1921)^(operation_194_1877));
            operation_194_1877 <= ((operation_194_1919)*(operation_194_5597));
            operation_194_1879 <= ((operation_194_1917)^(operation_194_1880));
            operation_194_1880 <= ((operation_194_1915)*(operation_194_5597));
            operation_194_1882 <= ((operation_194_1913)^(operation_194_1883));
            operation_194_1883 <= ((operation_194_1911)*(operation_194_5597));
            operation_194_1885 <= ((operation_194_1909)^(operation_194_1886));
            operation_194_1886 <= ((operation_194_1907)*(operation_194_5597));
            operation_194_1888 <= ((operation_194_1905)^(operation_194_1889));
            operation_194_1889 <= ((operation_194_1903)*(operation_194_5597));
            operation_194_1891 <= ((operation_194_1901)^(operation_194_1892));
            operation_194_1892 <= ((operation_194_1899)*(operation_194_5597));
            operation_194_1894 <= ((operation_194_77)^(operation_194_1898));
            operation_194_1896 <= ((operation_194_93)^(operation_194_1897));
            operation_194_1899 <= ((operation_194_1900)&(operation_194_5557));
            operation_194_1900 <= ((operation_194_1902)>>(operation_194_2119));
            operation_194_1901 <= ((operation_194_1902)<<(operation_194_5557));
            operation_194_1903 <= ((operation_194_1904)&(operation_194_5557));
            operation_194_1904 <= ((operation_194_1906)>>(operation_194_2119));
            operation_194_1905 <= ((operation_194_1906)<<(operation_194_5557));
            operation_194_1907 <= ((operation_194_1908)&(operation_194_5557));
            operation_194_1908 <= ((operation_194_1910)>>(operation_194_2119));
            operation_194_1909 <= ((operation_194_1910)<<(operation_194_5557));
            operation_194_1911 <= ((operation_194_1912)&(operation_194_5557));
            operation_194_1912 <= ((operation_194_1914)>>(operation_194_2119));
            operation_194_1913 <= ((operation_194_1914)<<(operation_194_5557));
            operation_194_1915 <= ((operation_194_1916)&(operation_194_5557));
            operation_194_1916 <= ((operation_194_1918)>>(operation_194_2119));
            operation_194_1917 <= ((operation_194_1918)<<(operation_194_5557));
            operation_194_1919 <= ((operation_194_1920)&(operation_194_5557));
            operation_194_1920 <= ((operation_194_1922)>>(operation_194_2119));
            operation_194_1921 <= ((operation_194_1922)<<(operation_194_5557));
            operation_194_1923 <= ((operation_194_1924)&(operation_194_5557));
            operation_194_1924 <= ((operation_194_1926)>>(operation_194_2119));
            operation_194_1925 <= ((operation_194_1926)<<(operation_194_5557));
            operation_194_1927 <= ((operation_194_1928)&(operation_194_5557));
            operation_194_1928 <= ((operation_194_1930)>>(operation_194_2119));
            operation_194_1929 <= ((operation_194_1930)<<(operation_194_5557));
            operation_194_1932 <= ((operation_194_1993)^(operation_194_1933));
            operation_194_1933 <= ((operation_194_1991)*(operation_194_5597));
            operation_194_1935 <= ((operation_194_1989)^(operation_194_1936));
            operation_194_1936 <= ((operation_194_1987)*(operation_194_5597));
            operation_194_1938 <= ((operation_194_1985)^(operation_194_1939));
            operation_194_1939 <= ((operation_194_1983)*(operation_194_5597));
            operation_194_1941 <= ((operation_194_1981)^(operation_194_1942));
            operation_194_1942 <= ((operation_194_1979)*(operation_194_5597));
            operation_194_1944 <= ((operation_194_1977)^(operation_194_1945));
            operation_194_1945 <= ((operation_194_1975)*(operation_194_5597));
            operation_194_1947 <= ((operation_194_1973)^(operation_194_1948));
            operation_194_1948 <= ((operation_194_1971)*(operation_194_5597));
            operation_194_1950 <= ((operation_194_1969)^(operation_194_1951));
            operation_194_1951 <= ((operation_194_1967)*(operation_194_5597));
            operation_194_1953 <= ((operation_194_1965)^(operation_194_1954));
            operation_194_1954 <= ((operation_194_1963)*(operation_194_5597));
            operation_194_1956 <= ((operation_194_5)^(operation_194_1960));
            operation_194_1958 <= ((operation_194_53)^(operation_194_1959));
            operation_194_1963 <= ((operation_194_1964)&(operation_194_5557));
            operation_194_1964 <= ((operation_194_1966)>>(operation_194_2119));
            operation_194_1965 <= ((operation_194_1966)<<(operation_194_5557));
            operation_194_1967 <= ((operation_194_1968)&(operation_194_5557));
            operation_194_1968 <= ((operation_194_1970)>>(operation_194_2119));
            operation_194_1969 <= ((operation_194_1970)<<(operation_194_5557));
            operation_194_1971 <= ((operation_194_1972)&(operation_194_5557));
            operation_194_1972 <= ((operation_194_1974)>>(operation_194_2119));
            operation_194_1973 <= ((operation_194_1974)<<(operation_194_5557));
            operation_194_1975 <= ((operation_194_1976)&(operation_194_5557));
            operation_194_1976 <= ((operation_194_1978)>>(operation_194_2119));
            operation_194_1977 <= ((operation_194_1978)<<(operation_194_5557));
            operation_194_1979 <= ((operation_194_1980)&(operation_194_5557));
            operation_194_1980 <= ((operation_194_1982)>>(operation_194_2119));
            operation_194_1981 <= ((operation_194_1982)<<(operation_194_5557));
            operation_194_1983 <= ((operation_194_1984)&(operation_194_5557));
            operation_194_1984 <= ((operation_194_1986)>>(operation_194_2119));
            operation_194_1985 <= ((operation_194_1986)<<(operation_194_5557));
            operation_194_1987 <= ((operation_194_1988)&(operation_194_5557));
            operation_194_1988 <= ((operation_194_1990)>>(operation_194_2119));
            operation_194_1989 <= ((operation_194_1990)<<(operation_194_5557));
            operation_194_1991 <= ((operation_194_1992)&(operation_194_5557));
            operation_194_1992 <= ((operation_194_1994)>>(operation_194_2119));
            operation_194_1993 <= ((operation_194_1994)<<(operation_194_5557));
            operation_194_1997 <= ((operation_194_2068)^(operation_194_2097));
            operation_194_2000 <= ((operation_194_2066)^(operation_194_2095));
            operation_194_2003 <= ((operation_194_2064)^(operation_194_2093));
            operation_194_2006 <= ((operation_194_2062)^(operation_194_2091));
            operation_194_2008 <= ((operation_194_2024)^(operation_194_2097));
            operation_194_2010 <= ((operation_194_2022)^(operation_194_2093));
            operation_194_2012 <= ((operation_194_2019)^(operation_194_5557));
            operation_194_2014 <= ((operation_194_45)^(operation_194_2018));
            operation_194_2016 <= ((operation_194_61)^(operation_194_2017));
            operation_194_2022 <= ((operation_194_2023)^(operation_194_2064));
            operation_194_2023 <= ((operation_194_2063)^(operation_194_2094));
            operation_194_2024 <= ((operation_194_2025)^(operation_194_2068));
            operation_194_2025 <= ((operation_194_2067)^(operation_194_2098));
            operation_194_2027 <= ((operation_194_2098)^(operation_194_2068));
            operation_194_2029 <= ((operation_194_2097)^(operation_194_2067));
            operation_194_2031 <= ((operation_194_2096)^(operation_194_2066));
            operation_194_2033 <= ((operation_194_2095)^(operation_194_2065));
            operation_194_2035 <= ((operation_194_2094)^(operation_194_2064));
            operation_194_2037 <= ((operation_194_2093)^(operation_194_2063));
            operation_194_2039 <= ((operation_194_2092)^(operation_194_2062));
            operation_194_2041 <= ((operation_194_2091)^(operation_194_2061));
            operation_194_2043 <= ((operation_194_2059)^(operation_194_2095));
            operation_194_2045 <= ((operation_194_2057)^(operation_194_2091));
            operation_194_2047 <= ((operation_194_21)^(operation_194_2054));
            operation_194_2057 <= ((operation_194_2058)^(operation_194_2062));
            operation_194_2058 <= ((operation_194_2061)^(operation_194_2092));
            operation_194_2059 <= ((operation_194_2060)^(operation_194_2066));
            operation_194_2060 <= ((operation_194_2065)^(operation_194_2096));
            operation_194_2072 <= ((operation_194_13)^(operation_194_2087));
            operation_194_2074 <= ((operation_194_29)^(operation_194_2085));
            operation_194_2089_latch <= (operation_194_2089);
            operation_194_2090_latch <= (operation_194_2090);
            operation_194_2099_latch <= (operation_194_2099);
            operation_194_2100_latch <= (operation_194_2100);
            operation_194_2101_latch <= (operation_194_2101);
            operation_194_2102_latch <= (operation_194_2102);
            operation_194_2103_latch <= (operation_194_2103);
            operation_194_2104_latch <= (operation_194_2104);
            operation_194_2105_latch <= (operation_194_2105);
            operation_194_2106_latch <= (operation_194_2106);
            operation_194_2107_latch <= (operation_194_2107);
            operation_194_2108_latch <= (operation_194_2108);
            operation_194_2109_latch <= (operation_194_2109);
            operation_194_2110_latch <= (operation_194_2110);
            operation_194_2111_latch <= (operation_194_2111);
            operation_194_2112_latch <= (operation_194_2112);
            operation_194_2113_latch <= (operation_194_2113);
            operation_194_2114_latch <= (operation_194_2114);
            operation_194_2115_latch <= (operation_194_2115);
            operation_194_2116_latch <= (operation_194_2116);
            operation_194_126 <= ((operation_194_123)^(operation_194_125));
            operation_194_6 <= ((operation_194_3)^(operation_194_5));
            operation_194_22 <= ((operation_194_19)^(operation_194_21));
            operation_194_38 <= ((operation_194_35)^(operation_194_37));
            operation_194_54 <= ((operation_194_51)^(operation_194_53));
            operation_194_70 <= ((operation_194_67)^(operation_194_69));
            operation_194_86 <= ((operation_194_83)^(operation_194_85));
            operation_194_102 <= ((operation_194_99)^(operation_194_101));
            operation_194_118 <= ((operation_194_115)^(operation_194_117));
            operation_194_14 <= ((operation_194_11)^(operation_194_13));
            operation_194_30 <= ((operation_194_27)^(operation_194_29));
            operation_194_46 <= ((operation_194_43)^(operation_194_45));
            operation_194_62 <= ((operation_194_59)^(operation_194_61));
            operation_194_78 <= ((operation_194_75)^(operation_194_77));
            operation_194_94 <= ((operation_194_91)^(operation_194_93));
            operation_194_110 <= ((operation_194_107)^(operation_194_109));
            control_194_follow <= (control_194_end);
            control_194_83 <= (control_194_82);
            control_194_82 <= (control_194_81);
            control_194_81 <= (control_194_80);
            control_194_80 <= (control_194_79);
            control_194_79 <= (control_194_78);
            control_194_78 <= (control_194_77);
            control_194_77 <= (control_194_76);
            control_194_76 <= (control_194_75);
            control_194_75 <= (control_194_74);
            control_194_74 <= (control_194_73);
            control_194_73 <= (control_194_72);
            control_194_72 <= (control_194_71);
            control_194_71 <= (control_194_70);
            control_194_70 <= (control_194_69);
            control_194_69 <= (control_194_68);
            control_194_68 <= (control_194_67);
            control_194_67 <= (control_194_66);
            control_194_66 <= (control_194_65);
            control_194_65 <= (control_194_64);
            control_194_64 <= (control_194_63);
            control_194_63 <= (control_194_62);
            control_194_62 <= (control_194_61);
            control_194_61 <= (control_194_60);
            control_194_60 <= (control_194_59);
            control_194_59 <= (control_194_58);
            control_194_58 <= (control_194_57);
            control_194_57 <= (control_194_56);
            control_194_56 <= (control_194_55);
            control_194_55 <= (control_194_54);
            control_194_54 <= (control_194_53);
            control_194_53 <= (control_194_52);
            control_194_52 <= (control_194_51);
            control_194_51 <= (control_194_50);
            control_194_50 <= (control_194_49);
            control_194_49 <= (control_194_48);
            control_194_48 <= (control_194_47);
            control_194_47 <= (control_194_46);
            control_194_46 <= (control_194_45);
            control_194_45 <= (control_194_44);
            control_194_44 <= (control_194_43);
            control_194_43 <= (control_194_42);
            control_194_42 <= (control_194_41);
            control_194_41 <= (control_194_40);
            control_194_40 <= (control_194_39);
            control_194_39 <= (control_194_38);
            control_194_38 <= (control_194_37);
            control_194_37 <= (control_194_36);
            control_194_36 <= (control_194_35);
            control_194_35 <= (control_194_34);
            control_194_34 <= (control_194_33);
            control_194_33 <= (control_194_32);
            control_194_32 <= (control_194_31);
            control_194_31 <= (control_194_30);
            control_194_30 <= (control_194_29);
            control_194_29 <= (control_194_28);
            control_194_28 <= (control_194_27);
            control_194_27 <= (control_194_26);
            control_194_26 <= (control_194_25);
            control_194_25 <= (control_194_24);
            control_194_24 <= (control_194_23);
            control_194_23 <= (control_194_22);
            control_194_22 <= (control_194_21);
            control_194_21 <= (control_194_20);
            control_194_20 <= (control_194_19);
            control_194_19 <= (control_194_18);
            control_194_18 <= (control_194_17);
            control_194_17 <= (control_194_16);
            control_194_16 <= (control_194_15);
            control_194_15 <= (control_194_14);
            control_194_14 <= (control_194_13);
            control_194_13 <= (control_194_12);
            control_194_12 <= (control_194_11);
            control_194_11 <= (control_194_10);
            control_194_10 <= (control_194_9);
            control_194_9 <= (control_194_8);
            control_194_8 <= (control_194_7);
            control_194_7 <= (control_194_6);
            control_194_6 <= (control_194_5);
            control_194_5 <= (control_194_4);
            control_194_4 <= (control_194_3);
            control_194_3 <= (control_194_2);
            control_194_2 <= (control_194_1);
            control_194_1 <= (control_194_start);
            input_key_194_follow <= (input_key_194);
            input_in_194_follow <= (input_in_194);
            lookup_sbox_0_output <= ((lookup_sbox_0_enable)?(sbox_0[(lookup_sbox_0_0)]):(lookup_sbox_0_output));
            lookup_sbox_1_output <= ((lookup_sbox_1_enable)?(sbox_1[(lookup_sbox_1_0)]):(lookup_sbox_1_output));
            lookup_sbox_2_output <= ((lookup_sbox_2_enable)?(sbox_2[(lookup_sbox_2_0)]):(lookup_sbox_2_output));
            lookup_sbox_3_output <= ((lookup_sbox_3_enable)?(sbox_3[(lookup_sbox_3_0)]):(lookup_sbox_3_output));
            lookup_sbox_4_output <= ((lookup_sbox_4_enable)?(sbox_4[(lookup_sbox_4_0)]):(lookup_sbox_4_output));
            lookup_sbox_5_output <= ((lookup_sbox_5_enable)?(sbox_5[(lookup_sbox_5_0)]):(lookup_sbox_5_output));
            lookup_sbox_6_output <= ((lookup_sbox_6_enable)?(sbox_6[(lookup_sbox_6_0)]):(lookup_sbox_6_output));
            lookup_sbox_7_output <= ((lookup_sbox_7_enable)?(sbox_7[(lookup_sbox_7_0)]):(lookup_sbox_7_output));
            lookup_sbox_8_output <= ((lookup_sbox_8_enable)?(sbox_8[(lookup_sbox_8_0)]):(lookup_sbox_8_output));
            lookup_sbox_9_output <= ((lookup_sbox_9_enable)?(sbox_9[(lookup_sbox_9_0)]):(lookup_sbox_9_output));
            lookup_sbox_10_output <= ((lookup_sbox_10_enable)?(sbox_10[(lookup_sbox_10_0)]):(lookup_sbox_10_output));
            lookup_sbox_11_output <= ((lookup_sbox_11_enable)?(sbox_11[(lookup_sbox_11_0)]):(lookup_sbox_11_output));
            lookup_sbox_12_output <= ((lookup_sbox_12_enable)?(sbox_12[(lookup_sbox_12_0)]):(lookup_sbox_12_output));
            lookup_sbox_13_output <= ((lookup_sbox_13_enable)?(sbox_13[(lookup_sbox_13_0)]):(lookup_sbox_13_output));
            lookup_sbox_14_output <= ((lookup_sbox_14_enable)?(sbox_14[(lookup_sbox_14_0)]):(lookup_sbox_14_output));
            lookup_sbox_15_output <= ((lookup_sbox_15_enable)?(sbox_15[(lookup_sbox_15_0)]):(lookup_sbox_15_output));
            lookup_sbox_16_output <= ((lookup_sbox_16_enable)?(sbox_16[(lookup_sbox_16_0)]):(lookup_sbox_16_output));
            lookup_sbox_17_output <= ((lookup_sbox_17_enable)?(sbox_17[(lookup_sbox_17_0)]):(lookup_sbox_17_output));
            lookup_sbox_18_output <= ((lookup_sbox_18_enable)?(sbox_18[(lookup_sbox_18_0)]):(lookup_sbox_18_output));
            lookup_sbox_19_output <= ((lookup_sbox_19_enable)?(sbox_19[(lookup_sbox_19_0)]):(lookup_sbox_19_output));
            lookup_sbox_20_output <= ((lookup_sbox_20_enable)?(sbox_20[(lookup_sbox_20_0)]):(lookup_sbox_20_output));
            lookup_sbox_21_output <= ((lookup_sbox_21_enable)?(sbox_21[(lookup_sbox_21_0)]):(lookup_sbox_21_output));
            lookup_sbox_22_output <= ((lookup_sbox_22_enable)?(sbox_22[(lookup_sbox_22_0)]):(lookup_sbox_22_output));
            lookup_sbox_23_output <= ((lookup_sbox_23_enable)?(sbox_23[(lookup_sbox_23_0)]):(lookup_sbox_23_output));
            lookup_sbox_24_output <= ((lookup_sbox_24_enable)?(sbox_24[(lookup_sbox_24_0)]):(lookup_sbox_24_output));
            lookup_sbox_25_output <= ((lookup_sbox_25_enable)?(sbox_25[(lookup_sbox_25_0)]):(lookup_sbox_25_output));
            lookup_sbox_26_output <= ((lookup_sbox_26_enable)?(sbox_26[(lookup_sbox_26_0)]):(lookup_sbox_26_output));
            lookup_sbox_27_output <= ((lookup_sbox_27_enable)?(sbox_27[(lookup_sbox_27_0)]):(lookup_sbox_27_output));
            lookup_sbox_28_output <= ((lookup_sbox_28_enable)?(sbox_28[(lookup_sbox_28_0)]):(lookup_sbox_28_output));
            lookup_sbox_29_output <= ((lookup_sbox_29_enable)?(sbox_29[(lookup_sbox_29_0)]):(lookup_sbox_29_output));
            lookup_sbox_30_output <= ((lookup_sbox_30_enable)?(sbox_30[(lookup_sbox_30_0)]):(lookup_sbox_30_output));
            lookup_sbox_31_output <= ((lookup_sbox_31_enable)?(sbox_31[(lookup_sbox_31_0)]):(lookup_sbox_31_output));
            startfollow <= (start);
        end
endmodule // end of module AES128_encrypt
