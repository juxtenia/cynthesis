module AES128_encrypt( input clk, input rst, input start, input [127:0] in, input [127:0] key, output reg finish, output reg [127:0] AES128_encrypt);
wire [127:0] return_274;
wire [7:0] operation_274_1665;
wire [7:0] operation_274_1689;
wire [7:0] operation_274_1673;
wire [7:0] operation_274_1633;
wire [7:0] operation_274_1681;
wire [7:0] operation_274_1657;
wire [7:0] operation_274_1641;
wire [7:0] operation_274_1601;
wire [7:0] operation_274_1649;
wire [7:0] operation_274_1625;
wire [7:0] operation_274_1609;
wire [7:0] operation_274_1569;
wire [7:0] operation_274_1617;
wire [7:0] operation_274_1593;
wire [7:0] operation_274_1577;
wire [7:0] operation_274_1585;
reg signed [31:0] operation_274_1664;
reg signed [31:0] operation_274_1688;
reg signed [31:0] operation_274_1672;
reg signed [31:0] operation_274_1632;
reg signed [31:0] operation_274_1680;
reg signed [31:0] operation_274_1656;
reg signed [31:0] operation_274_1640;
reg signed [31:0] operation_274_1600;
reg signed [31:0] operation_274_1648;
reg signed [31:0] operation_274_1624;
reg signed [31:0] operation_274_1608;
reg signed [31:0] operation_274_1568;
reg signed [31:0] operation_274_1616;
reg signed [31:0] operation_274_1592;
reg signed [31:0] operation_274_1576;
reg signed [31:0] operation_274_1584;
wire signed [31:0] operation_274_1685;
wire signed [31:0] operation_274_1669;
wire signed [31:0] operation_274_1653;
wire signed [31:0] operation_274_1637;
wire signed [31:0] operation_274_1621;
wire signed [31:0] operation_274_1605;
wire signed [31:0] operation_274_1589;
wire signed [31:0] operation_274_1573;
wire signed [31:0] operation_274_1565;
wire signed [31:0] operation_274_1581;
wire signed [31:0] operation_274_1597;
wire signed [31:0] operation_274_1613;
wire signed [31:0] operation_274_1629;
wire signed [31:0] operation_274_1645;
wire signed [31:0] operation_274_1661;
wire signed [31:0] operation_274_1677;
reg [7:0] operation_274_1338_latch;
wire [7:0] operation_274_1338;
reg [7:0] operation_274_1328_latch;
wire [7:0] operation_274_1328;
reg [7:0] operation_274_1318_latch;
wire [7:0] operation_274_1318;
reg [7:0] operation_274_1308_latch;
wire [7:0] operation_274_1308;
reg [7:0] operation_274_1298_latch;
wire [7:0] operation_274_1298;
reg [7:0] operation_274_1288_latch;
wire [7:0] operation_274_1288;
reg [7:0] operation_274_1278_latch;
wire [7:0] operation_274_1278;
reg [7:0] operation_274_1268_latch;
wire [7:0] operation_274_1268;
reg [7:0] operation_274_1273_latch;
wire [7:0] operation_274_1273;
reg [7:0] operation_274_1283_latch;
wire [7:0] operation_274_1283;
reg [7:0] operation_274_1293_latch;
wire [7:0] operation_274_1293;
reg [7:0] operation_274_1303_latch;
wire [7:0] operation_274_1303;
reg [7:0] operation_274_1313_latch;
wire [7:0] operation_274_1313;
reg [7:0] operation_274_1323_latch;
wire [7:0] operation_274_1323;
reg [7:0] operation_274_1333_latch;
wire [7:0] operation_274_1333;
reg [7:0] operation_274_1343_latch;
wire [7:0] operation_274_1343;
wire [7:0] operation_274_5146;
wire [7:0] operation_274_5145;
wire [7:0] operation_274_5144;
wire [7:0] operation_274_5143;
wire [7:0] operation_274_5142;
wire [7:0] operation_274_5141;
wire [7:0] operation_274_5140;
wire [7:0] operation_274_5139;
wire [7:0] operation_274_5138;
wire [7:0] operation_274_5137;
wire [7:0] operation_274_5136;
wire [7:0] operation_274_5135;
wire [7:0] operation_274_5134;
wire [7:0] operation_274_5133;
wire [7:0] operation_274_5132;
wire [7:0] operation_274_5131;
reg signed [31:0] operation_274_5162;
reg signed [31:0] operation_274_5161;
reg signed [31:0] operation_274_5160;
reg signed [31:0] operation_274_5159;
reg signed [31:0] operation_274_5158;
reg signed [31:0] operation_274_5157;
reg signed [31:0] operation_274_5156;
reg signed [31:0] operation_274_5155;
reg signed [31:0] operation_274_5154;
reg signed [31:0] operation_274_5153;
reg signed [31:0] operation_274_5152;
reg signed [31:0] operation_274_5151;
reg signed [31:0] operation_274_5150;
reg signed [31:0] operation_274_5149;
reg signed [31:0] operation_274_5148;
reg signed [31:0] operation_274_5147;
wire signed [31:0] operation_274_5180;
wire signed [31:0] operation_274_5179;
wire signed [31:0] operation_274_5178;
wire signed [31:0] operation_274_5177;
wire signed [31:0] operation_274_5176;
wire signed [31:0] operation_274_5175;
wire signed [31:0] operation_274_5174;
wire signed [31:0] operation_274_5173;
wire signed [31:0] operation_274_5171;
wire signed [31:0] operation_274_5170;
wire signed [31:0] operation_274_5169;
wire signed [31:0] operation_274_5168;
wire signed [31:0] operation_274_5167;
wire signed [31:0] operation_274_5166;
wire signed [31:0] operation_274_5165;
wire signed [31:0] operation_274_5163;
wire [7:0] operation_274_5197;
wire [7:0] operation_274_5196;
wire [7:0] operation_274_5195;
wire [7:0] operation_274_5194;
wire [7:0] operation_274_5193;
wire [7:0] operation_274_5192;
wire [7:0] operation_274_5191;
wire [7:0] operation_274_5190;
wire [7:0] operation_274_5189;
wire [7:0] operation_274_5188;
wire [7:0] operation_274_5187;
wire [7:0] operation_274_5186;
wire [7:0] operation_274_5185;
wire [7:0] operation_274_5184;
wire [7:0] operation_274_5183;
wire [7:0] operation_274_5182;
reg signed [31:0] operation_274_5214;
reg signed [31:0] operation_274_5213;
reg signed [31:0] operation_274_5212;
reg signed [31:0] operation_274_5211;
reg signed [31:0] operation_274_5210;
reg signed [31:0] operation_274_5209;
reg signed [31:0] operation_274_5208;
reg signed [31:0] operation_274_5207;
reg signed [31:0] operation_274_5206;
reg signed [31:0] operation_274_5205;
reg signed [31:0] operation_274_5204;
reg signed [31:0] operation_274_5203;
reg signed [31:0] operation_274_5202;
reg signed [31:0] operation_274_5201;
reg signed [31:0] operation_274_5200;
reg signed [31:0] operation_274_5199;
wire signed [31:0] operation_274_5232;
wire signed [31:0] operation_274_5231;
wire signed [31:0] operation_274_5230;
wire signed [31:0] operation_274_5229;
wire signed [31:0] operation_274_5228;
wire signed [31:0] operation_274_5227;
wire signed [31:0] operation_274_5226;
wire signed [31:0] operation_274_5225;
wire signed [31:0] operation_274_5224;
wire signed [31:0] operation_274_5223;
wire signed [31:0] operation_274_5222;
wire signed [31:0] operation_274_5221;
wire signed [31:0] operation_274_5220;
wire signed [31:0] operation_274_5219;
wire signed [31:0] operation_274_5218;
wire signed [31:0] operation_274_5217;
wire [7:0] operation_274_5252;
wire [7:0] operation_274_5251;
wire [7:0] operation_274_5250;
wire [7:0] operation_274_5249;
wire [7:0] operation_274_5248;
wire [7:0] operation_274_5247;
wire [7:0] operation_274_5246;
wire [7:0] operation_274_5245;
wire [7:0] operation_274_5244;
wire [7:0] operation_274_5243;
wire [7:0] operation_274_5242;
wire [7:0] operation_274_5241;
wire [7:0] operation_274_5240;
wire [7:0] operation_274_5239;
wire [7:0] operation_274_5238;
wire [7:0] operation_274_5237;
reg signed [31:0] operation_274_5272;
reg signed [31:0] operation_274_5271;
reg signed [31:0] operation_274_5270;
reg signed [31:0] operation_274_5269;
reg signed [31:0] operation_274_5268;
reg signed [31:0] operation_274_5267;
reg signed [31:0] operation_274_5266;
reg signed [31:0] operation_274_5265;
reg signed [31:0] operation_274_5264;
reg signed [31:0] operation_274_5263;
reg signed [31:0] operation_274_5262;
reg signed [31:0] operation_274_5261;
reg signed [31:0] operation_274_5260;
reg signed [31:0] operation_274_5259;
reg signed [31:0] operation_274_5258;
reg signed [31:0] operation_274_5257;
wire signed [31:0] operation_274_5292;
wire signed [31:0] operation_274_5291;
wire signed [31:0] operation_274_5290;
wire signed [31:0] operation_274_5289;
wire signed [31:0] operation_274_5288;
wire signed [31:0] operation_274_5287;
wire signed [31:0] operation_274_5286;
wire signed [31:0] operation_274_5285;
wire signed [31:0] operation_274_5284;
wire signed [31:0] operation_274_5283;
wire signed [31:0] operation_274_5282;
wire signed [31:0] operation_274_5281;
wire signed [31:0] operation_274_5280;
wire signed [31:0] operation_274_5279;
wire signed [31:0] operation_274_5278;
wire signed [31:0] operation_274_5277;
wire [7:0] operation_274_5312;
wire [7:0] operation_274_5311;
wire [7:0] operation_274_5310;
wire [7:0] operation_274_5309;
wire [7:0] operation_274_5308;
wire [7:0] operation_274_5307;
wire [7:0] operation_274_5306;
wire [7:0] operation_274_5305;
wire [7:0] operation_274_5304;
wire [7:0] operation_274_5303;
wire [7:0] operation_274_5302;
wire [7:0] operation_274_5301;
wire [7:0] operation_274_5300;
wire [7:0] operation_274_5299;
wire [7:0] operation_274_5298;
wire [7:0] operation_274_5297;
reg signed [31:0] operation_274_5332;
reg signed [31:0] operation_274_5331;
reg signed [31:0] operation_274_5330;
reg signed [31:0] operation_274_5329;
reg signed [31:0] operation_274_5328;
reg signed [31:0] operation_274_5327;
reg signed [31:0] operation_274_5326;
reg signed [31:0] operation_274_5325;
reg signed [31:0] operation_274_5324;
reg signed [31:0] operation_274_5323;
reg signed [31:0] operation_274_5322;
reg signed [31:0] operation_274_5321;
reg signed [31:0] operation_274_5320;
reg signed [31:0] operation_274_5319;
reg signed [31:0] operation_274_5318;
reg signed [31:0] operation_274_5317;
reg signed [31:0] operation_274_5352;
reg signed [31:0] operation_274_5351;
reg signed [31:0] operation_274_5350;
reg signed [31:0] operation_274_5349;
reg signed [31:0] operation_274_5348;
reg signed [31:0] operation_274_5347;
reg signed [31:0] operation_274_5346;
reg signed [31:0] operation_274_5345;
reg signed [31:0] operation_274_5344;
reg signed [31:0] operation_274_5343;
reg signed [31:0] operation_274_5342;
reg signed [31:0] operation_274_5341;
reg signed [31:0] operation_274_5340;
reg signed [31:0] operation_274_5339;
reg signed [31:0] operation_274_5338;
reg signed [31:0] operation_274_5337;
reg signed [31:0] operation_274_5376;
reg signed [31:0] operation_274_5375;
reg signed [31:0] operation_274_5374;
reg signed [31:0] operation_274_5373;
reg signed [31:0] operation_274_5372;
reg signed [31:0] operation_274_5371;
reg signed [31:0] operation_274_5370;
reg signed [31:0] operation_274_5369;
reg signed [31:0] operation_274_5368;
reg signed [31:0] operation_274_5367;
reg signed [31:0] operation_274_5366;
reg signed [31:0] operation_274_5365;
reg signed [31:0] operation_274_5364;
reg signed [31:0] operation_274_5363;
reg signed [31:0] operation_274_5362;
reg signed [31:0] operation_274_5361;
wire signed [31:0] operation_274_5360;
wire signed [31:0] operation_274_5359;
wire signed [31:0] operation_274_5358;
wire signed [31:0] operation_274_5357;
wire [7:0] operation_274_5416;
wire [7:0] operation_274_5415;
reg signed [31:0] operation_274_5414;
reg signed [31:0] operation_274_5413;
reg signed [31:0] operation_274_5412;
reg signed [31:0] operation_274_5411;
reg signed [31:0] operation_274_5410;
reg signed [31:0] operation_274_5409;
reg signed [31:0] operation_274_5408;
reg signed [31:0] operation_274_5407;
reg signed [31:0] operation_274_5406;
reg signed [31:0] operation_274_5405;
reg signed [31:0] operation_274_5404;
reg signed [31:0] operation_274_5403;
reg signed [31:0] operation_274_5402;
reg signed [31:0] operation_274_5401;
reg signed [31:0] operation_274_5400;
reg signed [31:0] operation_274_5399;
reg signed [31:0] operation_274_5398;
reg signed [31:0] operation_274_5397;
reg signed [31:0] operation_274_5396;
reg signed [31:0] operation_274_5395;
reg signed [31:0] operation_274_5394;
reg signed [31:0] operation_274_5393;
reg signed [31:0] operation_274_5392;
reg signed [31:0] operation_274_5391;
reg signed [31:0] operation_274_5390;
reg signed [31:0] operation_274_5389;
reg signed [31:0] operation_274_5388;
reg signed [31:0] operation_274_5387;
reg signed [31:0] operation_274_5386;
reg signed [31:0] operation_274_5385;
reg signed [31:0] operation_274_5384;
reg signed [31:0] operation_274_5383;
wire [7:0] operation_274_5382;
wire [7:0] operation_274_5381;
reg signed [31:0] operation_274_5440;
reg signed [31:0] operation_274_5439;
wire signed [31:0] operation_274_5438;
wire signed [31:0] operation_274_5437;
wire signed [31:0] operation_274_5436;
wire signed [31:0] operation_274_5435;
wire signed [31:0] operation_274_5434;
wire signed [31:0] operation_274_5433;
wire signed [31:0] operation_274_5432;
wire signed [31:0] operation_274_5431;
wire signed [31:0] operation_274_5430;
wire signed [31:0] operation_274_5429;
wire signed [31:0] operation_274_5428;
wire signed [31:0] operation_274_5427;
wire signed [31:0] operation_274_5426;
wire signed [31:0] operation_274_5425;
wire signed [31:0] operation_274_5424;
wire signed [31:0] operation_274_5423;
reg signed [31:0] operation_274_5422;
reg signed [31:0] operation_274_5421;
reg signed [31:0] operation_274_5464;
reg signed [31:0] operation_274_5463;
wire [7:0] operation_274_5462;
wire [7:0] operation_274_5461;
wire [7:0] operation_274_5460;
wire [7:0] operation_274_5459;
wire [7:0] operation_274_5458;
wire [7:0] operation_274_5457;
wire [7:0] operation_274_5456;
wire [7:0] operation_274_5455;
wire [7:0] operation_274_5454;
wire [7:0] operation_274_5453;
wire [7:0] operation_274_5452;
wire [7:0] operation_274_5451;
wire [7:0] operation_274_5450;
wire [7:0] operation_274_5449;
wire [7:0] operation_274_5448;
wire [7:0] operation_274_5447;
reg signed [31:0] operation_274_5446;
reg signed [31:0] operation_274_5445;
reg signed [31:0] operation_274_5485;
reg signed [31:0] operation_274_5484;
reg signed [31:0] operation_274_5483;
reg signed [31:0] operation_274_5482;
reg signed [31:0] operation_274_5481;
reg signed [31:0] operation_274_5480;
reg signed [31:0] operation_274_5479;
reg signed [31:0] operation_274_5478;
reg signed [31:0] operation_274_5477;
reg signed [31:0] operation_274_5476;
reg signed [31:0] operation_274_5475;
reg signed [31:0] operation_274_5474;
reg signed [31:0] operation_274_5473;
reg signed [31:0] operation_274_5472;
reg signed [31:0] operation_274_5471;
reg signed [31:0] operation_274_5470;
wire signed [31:0] operation_274_5507;
wire signed [31:0] operation_274_5506;
wire signed [31:0] operation_274_5505;
wire signed [31:0] operation_274_5504;
wire signed [31:0] operation_274_5503;
wire signed [31:0] operation_274_5502;
wire signed [31:0] operation_274_5501;
wire signed [31:0] operation_274_5500;
wire signed [31:0] operation_274_5499;
wire signed [31:0] operation_274_5498;
wire signed [31:0] operation_274_5497;
wire signed [31:0] operation_274_5496;
wire signed [31:0] operation_274_5495;
wire signed [31:0] operation_274_5494;
wire signed [31:0] operation_274_5493;
wire signed [31:0] operation_274_5492;
reg [7:0] operation_274_5536_latch;
wire [7:0] operation_274_5536;
reg [7:0] operation_274_5535_latch;
wire [7:0] operation_274_5535;
reg [7:0] operation_274_5534_latch;
wire [7:0] operation_274_5534;
reg [7:0] operation_274_5533_latch;
wire [7:0] operation_274_5533;
reg [7:0] operation_274_5532_latch;
wire [7:0] operation_274_5532;
reg [7:0] operation_274_5531_latch;
wire [7:0] operation_274_5531;
reg [7:0] operation_274_5530_latch;
wire [7:0] operation_274_5530;
reg [7:0] operation_274_5529_latch;
wire [7:0] operation_274_5529;
reg [7:0] operation_274_5528_latch;
wire [7:0] operation_274_5528;
reg [7:0] operation_274_5527_latch;
wire [7:0] operation_274_5527;
reg [7:0] operation_274_5526_latch;
wire [7:0] operation_274_5526;
reg [7:0] operation_274_5525_latch;
wire [7:0] operation_274_5525;
reg [7:0] operation_274_5524_latch;
wire [7:0] operation_274_5524;
reg [7:0] operation_274_5523_latch;
wire [7:0] operation_274_5523;
reg [7:0] operation_274_5522_latch;
wire [7:0] operation_274_5522;
reg [7:0] operation_274_5521_latch;
wire [7:0] operation_274_5521;
wire [7:0] operation_274_4717;
wire [7:0] operation_274_4716;
wire [7:0] operation_274_4715;
wire [7:0] operation_274_4714;
wire [7:0] operation_274_4713;
wire [7:0] operation_274_4712;
wire [7:0] operation_274_4711;
wire [7:0] operation_274_4710;
wire [7:0] operation_274_4709;
wire [7:0] operation_274_4708;
wire [7:0] operation_274_4707;
wire [7:0] operation_274_4706;
wire [7:0] operation_274_4705;
wire [7:0] operation_274_4704;
wire [7:0] operation_274_4703;
wire [7:0] operation_274_4702;
reg signed [31:0] operation_274_4733;
reg signed [31:0] operation_274_4732;
reg signed [31:0] operation_274_4731;
reg signed [31:0] operation_274_4730;
reg signed [31:0] operation_274_4729;
reg signed [31:0] operation_274_4728;
reg signed [31:0] operation_274_4727;
reg signed [31:0] operation_274_4726;
reg signed [31:0] operation_274_4725;
reg signed [31:0] operation_274_4724;
reg signed [31:0] operation_274_4723;
reg signed [31:0] operation_274_4722;
reg signed [31:0] operation_274_4721;
reg signed [31:0] operation_274_4720;
reg signed [31:0] operation_274_4719;
reg signed [31:0] operation_274_4718;
wire signed [31:0] operation_274_4751;
wire signed [31:0] operation_274_4750;
wire signed [31:0] operation_274_4749;
wire signed [31:0] operation_274_4748;
wire signed [31:0] operation_274_4747;
wire signed [31:0] operation_274_4746;
wire signed [31:0] operation_274_4745;
wire signed [31:0] operation_274_4744;
wire signed [31:0] operation_274_4742;
wire signed [31:0] operation_274_4741;
wire signed [31:0] operation_274_4740;
wire signed [31:0] operation_274_4739;
wire signed [31:0] operation_274_4738;
wire signed [31:0] operation_274_4737;
wire signed [31:0] operation_274_4736;
wire signed [31:0] operation_274_4734;
wire [7:0] operation_274_4768;
wire [7:0] operation_274_4767;
wire [7:0] operation_274_4766;
wire [7:0] operation_274_4765;
wire [7:0] operation_274_4764;
wire [7:0] operation_274_4763;
wire [7:0] operation_274_4762;
wire [7:0] operation_274_4761;
wire [7:0] operation_274_4760;
wire [7:0] operation_274_4759;
wire [7:0] operation_274_4758;
wire [7:0] operation_274_4757;
wire [7:0] operation_274_4756;
wire [7:0] operation_274_4755;
wire [7:0] operation_274_4754;
wire [7:0] operation_274_4753;
reg signed [31:0] operation_274_4785;
reg signed [31:0] operation_274_4784;
reg signed [31:0] operation_274_4783;
reg signed [31:0] operation_274_4782;
reg signed [31:0] operation_274_4781;
reg signed [31:0] operation_274_4780;
reg signed [31:0] operation_274_4779;
reg signed [31:0] operation_274_4778;
reg signed [31:0] operation_274_4777;
reg signed [31:0] operation_274_4776;
reg signed [31:0] operation_274_4775;
reg signed [31:0] operation_274_4774;
reg signed [31:0] operation_274_4773;
reg signed [31:0] operation_274_4772;
reg signed [31:0] operation_274_4771;
reg signed [31:0] operation_274_4770;
wire signed [31:0] operation_274_4803;
wire signed [31:0] operation_274_4802;
wire signed [31:0] operation_274_4801;
wire signed [31:0] operation_274_4800;
wire signed [31:0] operation_274_4799;
wire signed [31:0] operation_274_4798;
wire signed [31:0] operation_274_4797;
wire signed [31:0] operation_274_4796;
wire signed [31:0] operation_274_4795;
wire signed [31:0] operation_274_4794;
wire signed [31:0] operation_274_4793;
wire signed [31:0] operation_274_4792;
wire signed [31:0] operation_274_4791;
wire signed [31:0] operation_274_4790;
wire signed [31:0] operation_274_4789;
wire signed [31:0] operation_274_4788;
wire [7:0] operation_274_4823;
wire [7:0] operation_274_4822;
wire [7:0] operation_274_4821;
wire [7:0] operation_274_4820;
wire [7:0] operation_274_4819;
wire [7:0] operation_274_4818;
wire [7:0] operation_274_4817;
wire [7:0] operation_274_4816;
wire [7:0] operation_274_4815;
wire [7:0] operation_274_4814;
wire [7:0] operation_274_4813;
wire [7:0] operation_274_4812;
wire [7:0] operation_274_4811;
wire [7:0] operation_274_4810;
wire [7:0] operation_274_4809;
wire [7:0] operation_274_4808;
reg signed [31:0] operation_274_4843;
reg signed [31:0] operation_274_4842;
reg signed [31:0] operation_274_4841;
reg signed [31:0] operation_274_4840;
reg signed [31:0] operation_274_4839;
reg signed [31:0] operation_274_4838;
reg signed [31:0] operation_274_4837;
reg signed [31:0] operation_274_4836;
reg signed [31:0] operation_274_4835;
reg signed [31:0] operation_274_4834;
reg signed [31:0] operation_274_4833;
reg signed [31:0] operation_274_4832;
reg signed [31:0] operation_274_4831;
reg signed [31:0] operation_274_4830;
reg signed [31:0] operation_274_4829;
reg signed [31:0] operation_274_4828;
wire signed [31:0] operation_274_4863;
wire signed [31:0] operation_274_4862;
wire signed [31:0] operation_274_4861;
wire signed [31:0] operation_274_4860;
wire signed [31:0] operation_274_4859;
wire signed [31:0] operation_274_4858;
wire signed [31:0] operation_274_4857;
wire signed [31:0] operation_274_4856;
wire signed [31:0] operation_274_4855;
wire signed [31:0] operation_274_4854;
wire signed [31:0] operation_274_4853;
wire signed [31:0] operation_274_4852;
wire signed [31:0] operation_274_4851;
wire signed [31:0] operation_274_4850;
wire signed [31:0] operation_274_4849;
wire signed [31:0] operation_274_4848;
wire [7:0] operation_274_4883;
wire [7:0] operation_274_4882;
wire [7:0] operation_274_4881;
wire [7:0] operation_274_4880;
wire [7:0] operation_274_4879;
wire [7:0] operation_274_4878;
wire [7:0] operation_274_4877;
wire [7:0] operation_274_4876;
wire [7:0] operation_274_4875;
wire [7:0] operation_274_4874;
wire [7:0] operation_274_4873;
wire [7:0] operation_274_4872;
wire [7:0] operation_274_4871;
wire [7:0] operation_274_4870;
wire [7:0] operation_274_4869;
wire [7:0] operation_274_4868;
reg signed [31:0] operation_274_4903;
reg signed [31:0] operation_274_4902;
reg signed [31:0] operation_274_4901;
reg signed [31:0] operation_274_4900;
reg signed [31:0] operation_274_4899;
reg signed [31:0] operation_274_4898;
reg signed [31:0] operation_274_4897;
reg signed [31:0] operation_274_4896;
reg signed [31:0] operation_274_4895;
reg signed [31:0] operation_274_4894;
reg signed [31:0] operation_274_4893;
reg signed [31:0] operation_274_4892;
reg signed [31:0] operation_274_4891;
reg signed [31:0] operation_274_4890;
reg signed [31:0] operation_274_4889;
reg signed [31:0] operation_274_4888;
reg signed [31:0] operation_274_4923;
reg signed [31:0] operation_274_4922;
reg signed [31:0] operation_274_4921;
reg signed [31:0] operation_274_4920;
reg signed [31:0] operation_274_4919;
reg signed [31:0] operation_274_4918;
reg signed [31:0] operation_274_4917;
reg signed [31:0] operation_274_4916;
reg signed [31:0] operation_274_4915;
reg signed [31:0] operation_274_4914;
reg signed [31:0] operation_274_4913;
reg signed [31:0] operation_274_4912;
reg signed [31:0] operation_274_4911;
reg signed [31:0] operation_274_4910;
reg signed [31:0] operation_274_4909;
reg signed [31:0] operation_274_4908;
reg signed [31:0] operation_274_4947;
reg signed [31:0] operation_274_4946;
reg signed [31:0] operation_274_4945;
reg signed [31:0] operation_274_4944;
reg signed [31:0] operation_274_4943;
reg signed [31:0] operation_274_4942;
reg signed [31:0] operation_274_4941;
reg signed [31:0] operation_274_4940;
reg signed [31:0] operation_274_4939;
reg signed [31:0] operation_274_4938;
reg signed [31:0] operation_274_4937;
reg signed [31:0] operation_274_4936;
reg signed [31:0] operation_274_4935;
reg signed [31:0] operation_274_4934;
reg signed [31:0] operation_274_4933;
reg signed [31:0] operation_274_4932;
wire signed [31:0] operation_274_4931;
wire signed [31:0] operation_274_4930;
wire signed [31:0] operation_274_4929;
wire signed [31:0] operation_274_4928;
wire [7:0] operation_274_4987;
wire [7:0] operation_274_4986;
reg signed [31:0] operation_274_4985;
reg signed [31:0] operation_274_4984;
reg signed [31:0] operation_274_4983;
reg signed [31:0] operation_274_4982;
reg signed [31:0] operation_274_4981;
reg signed [31:0] operation_274_4980;
reg signed [31:0] operation_274_4979;
reg signed [31:0] operation_274_4978;
reg signed [31:0] operation_274_4977;
reg signed [31:0] operation_274_4976;
reg signed [31:0] operation_274_4975;
reg signed [31:0] operation_274_4974;
reg signed [31:0] operation_274_4973;
reg signed [31:0] operation_274_4972;
reg signed [31:0] operation_274_4971;
reg signed [31:0] operation_274_4970;
reg signed [31:0] operation_274_4969;
reg signed [31:0] operation_274_4968;
reg signed [31:0] operation_274_4967;
reg signed [31:0] operation_274_4966;
reg signed [31:0] operation_274_4965;
reg signed [31:0] operation_274_4964;
reg signed [31:0] operation_274_4963;
reg signed [31:0] operation_274_4962;
reg signed [31:0] operation_274_4961;
reg signed [31:0] operation_274_4960;
reg signed [31:0] operation_274_4959;
reg signed [31:0] operation_274_4958;
reg signed [31:0] operation_274_4957;
reg signed [31:0] operation_274_4956;
reg signed [31:0] operation_274_4955;
reg signed [31:0] operation_274_4954;
wire [7:0] operation_274_4953;
wire [7:0] operation_274_4952;
reg signed [31:0] operation_274_5011;
reg signed [31:0] operation_274_5010;
wire signed [31:0] operation_274_5009;
wire signed [31:0] operation_274_5008;
wire signed [31:0] operation_274_5007;
wire signed [31:0] operation_274_5006;
wire signed [31:0] operation_274_5005;
wire signed [31:0] operation_274_5004;
wire signed [31:0] operation_274_5003;
wire signed [31:0] operation_274_5002;
wire signed [31:0] operation_274_5001;
wire signed [31:0] operation_274_5000;
wire signed [31:0] operation_274_4999;
wire signed [31:0] operation_274_4998;
wire signed [31:0] operation_274_4997;
wire signed [31:0] operation_274_4996;
wire signed [31:0] operation_274_4995;
wire signed [31:0] operation_274_4994;
reg signed [31:0] operation_274_4993;
reg signed [31:0] operation_274_4992;
reg signed [31:0] operation_274_5035;
reg signed [31:0] operation_274_5034;
wire [7:0] operation_274_5033;
wire [7:0] operation_274_5032;
wire [7:0] operation_274_5031;
wire [7:0] operation_274_5030;
wire [7:0] operation_274_5029;
wire [7:0] operation_274_5028;
wire [7:0] operation_274_5027;
wire [7:0] operation_274_5026;
wire [7:0] operation_274_5025;
wire [7:0] operation_274_5024;
wire [7:0] operation_274_5023;
wire [7:0] operation_274_5022;
wire [7:0] operation_274_5021;
wire [7:0] operation_274_5020;
wire [7:0] operation_274_5019;
wire [7:0] operation_274_5018;
reg signed [31:0] operation_274_5017;
reg signed [31:0] operation_274_5016;
wire signed [31:0] operation_274_1663;
wire signed [31:0] operation_274_1687;
reg signed [31:0] operation_274_5056;
reg signed [31:0] operation_274_5055;
reg signed [31:0] operation_274_5054;
reg signed [31:0] operation_274_5053;
reg signed [31:0] operation_274_5052;
reg signed [31:0] operation_274_5051;
reg signed [31:0] operation_274_5050;
reg signed [31:0] operation_274_5049;
reg signed [31:0] operation_274_5048;
reg signed [31:0] operation_274_5047;
reg signed [31:0] operation_274_5046;
reg signed [31:0] operation_274_5045;
reg signed [31:0] operation_274_5044;
reg signed [31:0] operation_274_5043;
reg signed [31:0] operation_274_5042;
reg signed [31:0] operation_274_5041;
wire [7:0] operation_274_1537;
wire [7:0] operation_274_1561;
wire signed [31:0] operation_274_5078;
wire signed [31:0] operation_274_5077;
wire signed [31:0] operation_274_5076;
wire signed [31:0] operation_274_5075;
wire signed [31:0] operation_274_5074;
wire signed [31:0] operation_274_5073;
wire signed [31:0] operation_274_5072;
wire signed [31:0] operation_274_5071;
wire signed [31:0] operation_274_5070;
wire signed [31:0] operation_274_5069;
wire signed [31:0] operation_274_5068;
wire signed [31:0] operation_274_5067;
wire signed [31:0] operation_274_5066;
wire signed [31:0] operation_274_5065;
wire signed [31:0] operation_274_5064;
wire signed [31:0] operation_274_5063;
reg signed [31:0] operation_274_1536;
reg signed [31:0] operation_274_1560;
reg [7:0] operation_274_5107_latch;
wire [7:0] operation_274_5107;
reg [7:0] operation_274_5106_latch;
wire [7:0] operation_274_5106;
reg [7:0] operation_274_5105_latch;
wire [7:0] operation_274_5105;
reg [7:0] operation_274_5104_latch;
wire [7:0] operation_274_5104;
reg [7:0] operation_274_5103_latch;
wire [7:0] operation_274_5103;
reg [7:0] operation_274_5102_latch;
wire [7:0] operation_274_5102;
reg [7:0] operation_274_5101_latch;
wire [7:0] operation_274_5101;
reg [7:0] operation_274_5100_latch;
wire [7:0] operation_274_5100;
reg [7:0] operation_274_5099_latch;
wire [7:0] operation_274_5099;
reg [7:0] operation_274_5098_latch;
wire [7:0] operation_274_5098;
reg [7:0] operation_274_5097_latch;
wire [7:0] operation_274_5097;
reg [7:0] operation_274_5096_latch;
wire [7:0] operation_274_5096;
reg [7:0] operation_274_5095_latch;
wire [7:0] operation_274_5095;
reg [7:0] operation_274_5094_latch;
wire [7:0] operation_274_5094;
reg [7:0] operation_274_5093_latch;
wire [7:0] operation_274_5093;
reg [7:0] operation_274_5092_latch;
wire [7:0] operation_274_5092;
wire signed [31:0] operation_274_1671;
wire signed [31:0] operation_274_1535;
wire signed [31:0] operation_274_1679;
wire signed [31:0] operation_274_1655;
wire [7:0] operation_274_4288;
wire [7:0] operation_274_4287;
wire [7:0] operation_274_4286;
wire [7:0] operation_274_4285;
wire [7:0] operation_274_4284;
wire [7:0] operation_274_4283;
wire [7:0] operation_274_4282;
wire [7:0] operation_274_4281;
wire [7:0] operation_274_4280;
wire [7:0] operation_274_4279;
wire [7:0] operation_274_4278;
wire [7:0] operation_274_4277;
wire [7:0] operation_274_4276;
wire [7:0] operation_274_4275;
wire [7:0] operation_274_4274;
wire [7:0] operation_274_4273;
wire [7:0] operation_274_1545;
wire [7:0] operation_274_1505;
wire [7:0] operation_274_1553;
wire [7:0] operation_274_1529;
reg signed [31:0] operation_274_4304;
reg signed [31:0] operation_274_4303;
reg signed [31:0] operation_274_4302;
reg signed [31:0] operation_274_4301;
reg signed [31:0] operation_274_4300;
reg signed [31:0] operation_274_4299;
reg signed [31:0] operation_274_4298;
reg signed [31:0] operation_274_4297;
reg signed [31:0] operation_274_4296;
reg signed [31:0] operation_274_4295;
reg signed [31:0] operation_274_4294;
reg signed [31:0] operation_274_4293;
reg signed [31:0] operation_274_4292;
reg signed [31:0] operation_274_4291;
reg signed [31:0] operation_274_4290;
reg signed [31:0] operation_274_4289;
reg signed [31:0] operation_274_1544;
reg signed [31:0] operation_274_1504;
reg signed [31:0] operation_274_1552;
reg signed [31:0] operation_274_1528;
wire signed [31:0] operation_274_4322;
wire signed [31:0] operation_274_4321;
wire signed [31:0] operation_274_4320;
wire signed [31:0] operation_274_4319;
wire signed [31:0] operation_274_4318;
wire signed [31:0] operation_274_4317;
wire signed [31:0] operation_274_4316;
wire signed [31:0] operation_274_4315;
wire signed [31:0] operation_274_4313;
wire signed [31:0] operation_274_4312;
wire signed [31:0] operation_274_4311;
wire signed [31:0] operation_274_4310;
wire signed [31:0] operation_274_4309;
wire signed [31:0] operation_274_4308;
wire signed [31:0] operation_274_4307;
wire signed [31:0] operation_274_4305;
wire signed [31:0] operation_274_1639;
wire signed [31:0] operation_274_1503;
wire signed [31:0] operation_274_1551;
wire signed [31:0] operation_274_1623;
wire [7:0] operation_274_4339;
wire [7:0] operation_274_4338;
wire [7:0] operation_274_4337;
wire [7:0] operation_274_4336;
wire [7:0] operation_274_4335;
wire [7:0] operation_274_4334;
wire [7:0] operation_274_4333;
wire [7:0] operation_274_4332;
wire [7:0] operation_274_4331;
wire [7:0] operation_274_4330;
wire [7:0] operation_274_4329;
wire [7:0] operation_274_4328;
wire [7:0] operation_274_4327;
wire [7:0] operation_274_4326;
wire [7:0] operation_274_4325;
wire [7:0] operation_274_4324;
wire [7:0] operation_274_1513;
wire [7:0] operation_274_1473;
wire [7:0] operation_274_1521;
wire [7:0] operation_274_1497;
reg signed [31:0] operation_274_4356;
reg signed [31:0] operation_274_4355;
reg signed [31:0] operation_274_4354;
reg signed [31:0] operation_274_4353;
reg signed [31:0] operation_274_4352;
reg signed [31:0] operation_274_4351;
reg signed [31:0] operation_274_4350;
reg signed [31:0] operation_274_4349;
reg signed [31:0] operation_274_4348;
reg signed [31:0] operation_274_4347;
reg signed [31:0] operation_274_4346;
reg signed [31:0] operation_274_4345;
reg signed [31:0] operation_274_4344;
reg signed [31:0] operation_274_4343;
reg signed [31:0] operation_274_4342;
reg signed [31:0] operation_274_4341;
reg signed [31:0] operation_274_1512;
reg signed [31:0] operation_274_1472;
reg signed [31:0] operation_274_1520;
reg signed [31:0] operation_274_1496;
wire signed [31:0] operation_274_4374;
wire signed [31:0] operation_274_4373;
wire signed [31:0] operation_274_4372;
wire signed [31:0] operation_274_4371;
wire signed [31:0] operation_274_4370;
wire signed [31:0] operation_274_4369;
wire signed [31:0] operation_274_4368;
wire signed [31:0] operation_274_4367;
wire signed [31:0] operation_274_4366;
wire signed [31:0] operation_274_4365;
wire signed [31:0] operation_274_4364;
wire signed [31:0] operation_274_4363;
wire signed [31:0] operation_274_4362;
wire signed [31:0] operation_274_4361;
wire signed [31:0] operation_274_4360;
wire signed [31:0] operation_274_4359;
wire signed [31:0] operation_274_1607;
wire signed [31:0] operation_274_1471;
wire signed [31:0] operation_274_1519;
wire signed [31:0] operation_274_1591;
wire [7:0] operation_274_4394;
wire [7:0] operation_274_4393;
wire [7:0] operation_274_4392;
wire [7:0] operation_274_4391;
wire [7:0] operation_274_4390;
wire [7:0] operation_274_4389;
wire [7:0] operation_274_4388;
wire [7:0] operation_274_4387;
wire [7:0] operation_274_4386;
wire [7:0] operation_274_4385;
wire [7:0] operation_274_4384;
wire [7:0] operation_274_4383;
wire [7:0] operation_274_4382;
wire [7:0] operation_274_4381;
wire [7:0] operation_274_4380;
wire [7:0] operation_274_4379;
wire [7:0] operation_274_1481;
wire [7:0] operation_274_1441;
wire [7:0] operation_274_1489;
wire [7:0] operation_274_1465;
reg signed [31:0] operation_274_4414;
reg signed [31:0] operation_274_4413;
reg signed [31:0] operation_274_4412;
reg signed [31:0] operation_274_4411;
reg signed [31:0] operation_274_4410;
reg signed [31:0] operation_274_4409;
reg signed [31:0] operation_274_4408;
reg signed [31:0] operation_274_4407;
reg signed [31:0] operation_274_4406;
reg signed [31:0] operation_274_4405;
reg signed [31:0] operation_274_4404;
reg signed [31:0] operation_274_4403;
reg signed [31:0] operation_274_4402;
reg signed [31:0] operation_274_4401;
reg signed [31:0] operation_274_4400;
reg signed [31:0] operation_274_4399;
reg signed [31:0] operation_274_1480;
reg signed [31:0] operation_274_1440;
reg signed [31:0] operation_274_1488;
reg signed [31:0] operation_274_1464;
wire signed [31:0] operation_274_4434;
wire signed [31:0] operation_274_4433;
wire signed [31:0] operation_274_4432;
wire signed [31:0] operation_274_4431;
wire signed [31:0] operation_274_4430;
wire signed [31:0] operation_274_4429;
wire signed [31:0] operation_274_4428;
wire signed [31:0] operation_274_4427;
wire signed [31:0] operation_274_4426;
wire signed [31:0] operation_274_4425;
wire signed [31:0] operation_274_4424;
wire signed [31:0] operation_274_4423;
wire signed [31:0] operation_274_4422;
wire signed [31:0] operation_274_4421;
wire signed [31:0] operation_274_4420;
wire signed [31:0] operation_274_4419;
wire signed [31:0] operation_274_1575;
wire signed [31:0] operation_274_1439;
wire signed [31:0] operation_274_1487;
wire signed [31:0] operation_274_1463;
wire [7:0] operation_274_4454;
wire [7:0] operation_274_4453;
wire [7:0] operation_274_4452;
wire [7:0] operation_274_4451;
wire [7:0] operation_274_4450;
wire [7:0] operation_274_4449;
wire [7:0] operation_274_4448;
wire [7:0] operation_274_4447;
wire [7:0] operation_274_4446;
wire [7:0] operation_274_4445;
wire [7:0] operation_274_4444;
wire [7:0] operation_274_4443;
wire [7:0] operation_274_4442;
wire [7:0] operation_274_4441;
wire [7:0] operation_274_4440;
wire [7:0] operation_274_4439;
wire signed [31:0] operation_274_5164;
wire [7:0] operation_274_1449;
wire [7:0] operation_274_1433;
wire [7:0] operation_274_1457;
reg [7:0] operation_274_1423_latch;
wire [7:0] operation_274_1423;
reg signed [31:0] operation_274_4474;
reg signed [31:0] operation_274_4473;
reg signed [31:0] operation_274_4472;
reg signed [31:0] operation_274_4471;
reg signed [31:0] operation_274_4470;
reg signed [31:0] operation_274_4469;
reg signed [31:0] operation_274_4468;
reg signed [31:0] operation_274_4467;
reg signed [31:0] operation_274_4466;
reg signed [31:0] operation_274_4465;
reg signed [31:0] operation_274_4464;
reg signed [31:0] operation_274_4463;
reg signed [31:0] operation_274_4462;
reg signed [31:0] operation_274_4461;
reg signed [31:0] operation_274_4460;
reg signed [31:0] operation_274_4459;
wire [7:0] operation_274_5181;
reg signed [31:0] operation_274_1448;
reg signed [31:0] operation_274_1432;
reg signed [31:0] operation_274_1456;
reg signed [31:0] operation_274_4494;
reg signed [31:0] operation_274_4493;
reg signed [31:0] operation_274_4492;
reg signed [31:0] operation_274_4491;
reg signed [31:0] operation_274_4490;
reg signed [31:0] operation_274_4489;
reg signed [31:0] operation_274_4488;
reg signed [31:0] operation_274_4487;
reg signed [31:0] operation_274_4486;
reg signed [31:0] operation_274_4485;
reg signed [31:0] operation_274_4484;
reg signed [31:0] operation_274_4483;
reg signed [31:0] operation_274_4482;
reg signed [31:0] operation_274_4481;
reg signed [31:0] operation_274_4480;
reg signed [31:0] operation_274_4479;
reg signed [31:0] operation_274_5198;
wire signed [31:0] operation_274_1447;
wire signed [31:0] operation_274_1428;
wire signed [31:0] operation_274_1455;
reg signed [31:0] operation_274_4518;
reg signed [31:0] operation_274_4517;
reg signed [31:0] operation_274_4516;
reg signed [31:0] operation_274_4515;
reg signed [31:0] operation_274_4514;
reg signed [31:0] operation_274_4513;
reg signed [31:0] operation_274_4512;
reg signed [31:0] operation_274_4511;
reg signed [31:0] operation_274_4510;
reg signed [31:0] operation_274_4509;
reg signed [31:0] operation_274_4508;
reg signed [31:0] operation_274_4507;
reg signed [31:0] operation_274_4506;
reg signed [31:0] operation_274_4505;
reg signed [31:0] operation_274_4504;
reg signed [31:0] operation_274_4503;
wire signed [31:0] operation_274_4502;
wire signed [31:0] operation_274_4501;
wire signed [31:0] operation_274_4500;
wire signed [31:0] operation_274_4499;
wire signed [31:0] operation_274_5234;
wire signed [31:0] operation_274_5233;
wire signed [31:0] operation_274_5216;
wire signed [31:0] operation_274_5215;
reg [7:0] operation_274_1418_latch;
wire [7:0] operation_274_1418;
reg [7:0] operation_274_1408_latch;
wire [7:0] operation_274_1408;
reg [7:0] operation_274_1413_latch;
wire [7:0] operation_274_1413;
wire [7:0] operation_274_4558;
wire [7:0] operation_274_4557;
reg signed [31:0] operation_274_4556;
reg signed [31:0] operation_274_4555;
reg signed [31:0] operation_274_4554;
reg signed [31:0] operation_274_4553;
reg signed [31:0] operation_274_4552;
reg signed [31:0] operation_274_4551;
reg signed [31:0] operation_274_4550;
reg signed [31:0] operation_274_4549;
reg signed [31:0] operation_274_4548;
reg signed [31:0] operation_274_4547;
reg signed [31:0] operation_274_4546;
reg signed [31:0] operation_274_4545;
reg signed [31:0] operation_274_4544;
reg signed [31:0] operation_274_4543;
reg signed [31:0] operation_274_4542;
reg signed [31:0] operation_274_4541;
reg signed [31:0] operation_274_4540;
reg signed [31:0] operation_274_4539;
reg signed [31:0] operation_274_4538;
reg signed [31:0] operation_274_4537;
reg signed [31:0] operation_274_4536;
reg signed [31:0] operation_274_4535;
reg signed [31:0] operation_274_4534;
reg signed [31:0] operation_274_4533;
reg signed [31:0] operation_274_4532;
reg signed [31:0] operation_274_4531;
reg signed [31:0] operation_274_4530;
reg signed [31:0] operation_274_4529;
reg signed [31:0] operation_274_4528;
reg signed [31:0] operation_274_4527;
reg signed [31:0] operation_274_4526;
reg signed [31:0] operation_274_4525;
wire [7:0] operation_274_4524;
wire [7:0] operation_274_4523;
wire [7:0] operation_274_5254;
wire [7:0] operation_274_5253;
wire [7:0] operation_274_5236;
wire [7:0] operation_274_5235;
reg signed [31:0] operation_274_4582;
reg signed [31:0] operation_274_4581;
wire signed [31:0] operation_274_4580;
wire signed [31:0] operation_274_4579;
wire signed [31:0] operation_274_4578;
wire signed [31:0] operation_274_4577;
wire signed [31:0] operation_274_4576;
wire signed [31:0] operation_274_4575;
wire signed [31:0] operation_274_4574;
wire signed [31:0] operation_274_4573;
wire signed [31:0] operation_274_4572;
wire signed [31:0] operation_274_4571;
wire signed [31:0] operation_274_4570;
wire signed [31:0] operation_274_4569;
wire signed [31:0] operation_274_4568;
wire signed [31:0] operation_274_4567;
wire signed [31:0] operation_274_4566;
wire signed [31:0] operation_274_4565;
reg signed [31:0] operation_274_4564;
reg signed [31:0] operation_274_4563;
reg signed [31:0] operation_274_5274;
reg signed [31:0] operation_274_5273;
reg signed [31:0] operation_274_5256;
reg signed [31:0] operation_274_5255;
reg signed [31:0] operation_274_4606;
reg signed [31:0] operation_274_4605;
wire [7:0] operation_274_4604;
wire [7:0] operation_274_4603;
wire [7:0] operation_274_4602;
wire [7:0] operation_274_4601;
wire [7:0] operation_274_4600;
wire [7:0] operation_274_4599;
wire [7:0] operation_274_4598;
wire [7:0] operation_274_4597;
wire [7:0] operation_274_4596;
wire [7:0] operation_274_4595;
wire [7:0] operation_274_4594;
wire [7:0] operation_274_4593;
wire [7:0] operation_274_4592;
wire [7:0] operation_274_4591;
wire [7:0] operation_274_4590;
wire [7:0] operation_274_4589;
reg signed [31:0] operation_274_4588;
reg signed [31:0] operation_274_4587;
wire signed [31:0] operation_274_5294;
wire signed [31:0] operation_274_5293;
wire signed [31:0] operation_274_5276;
wire signed [31:0] operation_274_5275;
reg signed [31:0] operation_274_4627;
reg signed [31:0] operation_274_4626;
reg signed [31:0] operation_274_4625;
reg signed [31:0] operation_274_4624;
reg signed [31:0] operation_274_4623;
reg signed [31:0] operation_274_4622;
reg signed [31:0] operation_274_4621;
reg signed [31:0] operation_274_4620;
reg signed [31:0] operation_274_4619;
reg signed [31:0] operation_274_4618;
reg signed [31:0] operation_274_4617;
reg signed [31:0] operation_274_4616;
reg signed [31:0] operation_274_4615;
reg signed [31:0] operation_274_4614;
reg signed [31:0] operation_274_4613;
reg signed [31:0] operation_274_4612;
wire [7:0] operation_274_5314;
wire [7:0] operation_274_5313;
wire [7:0] operation_274_5296;
wire [7:0] operation_274_5295;
wire signed [31:0] operation_274_4649;
wire signed [31:0] operation_274_4648;
wire signed [31:0] operation_274_4647;
wire signed [31:0] operation_274_4646;
wire signed [31:0] operation_274_4645;
wire signed [31:0] operation_274_4644;
wire signed [31:0] operation_274_4643;
wire signed [31:0] operation_274_4642;
wire signed [31:0] operation_274_4641;
wire signed [31:0] operation_274_4640;
wire signed [31:0] operation_274_4639;
wire signed [31:0] operation_274_4638;
wire signed [31:0] operation_274_4637;
wire signed [31:0] operation_274_4636;
wire signed [31:0] operation_274_4635;
wire signed [31:0] operation_274_4634;
reg signed [31:0] operation_274_5334;
reg signed [31:0] operation_274_5333;
reg signed [31:0] operation_274_5316;
reg signed [31:0] operation_274_5315;
reg [7:0] operation_274_4678_latch;
wire [7:0] operation_274_4678;
reg [7:0] operation_274_4677_latch;
wire [7:0] operation_274_4677;
reg [7:0] operation_274_4676_latch;
wire [7:0] operation_274_4676;
reg [7:0] operation_274_4675_latch;
wire [7:0] operation_274_4675;
reg [7:0] operation_274_4674_latch;
wire [7:0] operation_274_4674;
reg [7:0] operation_274_4673_latch;
wire [7:0] operation_274_4673;
reg [7:0] operation_274_4672_latch;
wire [7:0] operation_274_4672;
reg [7:0] operation_274_4671_latch;
wire [7:0] operation_274_4671;
reg [7:0] operation_274_4670_latch;
wire [7:0] operation_274_4670;
reg [7:0] operation_274_4669_latch;
wire [7:0] operation_274_4669;
reg [7:0] operation_274_4668_latch;
wire [7:0] operation_274_4668;
reg [7:0] operation_274_4667_latch;
wire [7:0] operation_274_4667;
reg [7:0] operation_274_4666_latch;
wire [7:0] operation_274_4666;
reg [7:0] operation_274_4665_latch;
wire [7:0] operation_274_4665;
reg [7:0] operation_274_4664_latch;
wire [7:0] operation_274_4664;
reg [7:0] operation_274_4663_latch;
wire [7:0] operation_274_4663;
wire signed [31:0] operation_274_5354;
wire signed [31:0] operation_274_5353;
wire signed [31:0] operation_274_5336;
wire signed [31:0] operation_274_5335;
wire [7:0] operation_274_3859;
wire [7:0] operation_274_3858;
wire [7:0] operation_274_3857;
wire [7:0] operation_274_3856;
wire [7:0] operation_274_3855;
wire [7:0] operation_274_3854;
wire [7:0] operation_274_3853;
wire [7:0] operation_274_3852;
wire [7:0] operation_274_3851;
wire [7:0] operation_274_3850;
wire [7:0] operation_274_3849;
wire [7:0] operation_274_3848;
wire [7:0] operation_274_3847;
wire [7:0] operation_274_3846;
wire [7:0] operation_274_3845;
wire [7:0] operation_274_3844;
wire [7:0] operation_274_5378;
wire [7:0] operation_274_5377;
wire [7:0] operation_274_5356;
wire [7:0] operation_274_5355;
reg signed [31:0] operation_274_3875;
reg signed [31:0] operation_274_3874;
reg signed [31:0] operation_274_3873;
reg signed [31:0] operation_274_3872;
reg signed [31:0] operation_274_3871;
reg signed [31:0] operation_274_3870;
reg signed [31:0] operation_274_3869;
reg signed [31:0] operation_274_3868;
reg signed [31:0] operation_274_3867;
reg signed [31:0] operation_274_3866;
reg signed [31:0] operation_274_3865;
reg signed [31:0] operation_274_3864;
reg signed [31:0] operation_274_3863;
reg signed [31:0] operation_274_3862;
reg signed [31:0] operation_274_3861;
reg signed [31:0] operation_274_3860;
reg signed [31:0] operation_274_5418;
reg signed [31:0] operation_274_5417;
reg signed [31:0] operation_274_5380;
reg signed [31:0] operation_274_5379;
wire signed [31:0] operation_274_3893;
wire signed [31:0] operation_274_3892;
wire signed [31:0] operation_274_3891;
wire signed [31:0] operation_274_3890;
wire signed [31:0] operation_274_3889;
wire signed [31:0] operation_274_3888;
wire signed [31:0] operation_274_3887;
wire signed [31:0] operation_274_3886;
wire signed [31:0] operation_274_3884;
wire signed [31:0] operation_274_3883;
wire signed [31:0] operation_274_3882;
wire signed [31:0] operation_274_3881;
wire signed [31:0] operation_274_3880;
wire signed [31:0] operation_274_3879;
wire signed [31:0] operation_274_3878;
wire signed [31:0] operation_274_3876;
wire signed [31:0] operation_274_5442;
wire signed [31:0] operation_274_5441;
wire signed [31:0] operation_274_5420;
wire signed [31:0] operation_274_5419;
wire [7:0] operation_274_3910;
wire [7:0] operation_274_3909;
wire [7:0] operation_274_3908;
wire [7:0] operation_274_3907;
wire [7:0] operation_274_3906;
wire [7:0] operation_274_3905;
wire [7:0] operation_274_3904;
wire [7:0] operation_274_3903;
wire [7:0] operation_274_3902;
wire [7:0] operation_274_3901;
wire [7:0] operation_274_3900;
wire [7:0] operation_274_3899;
wire [7:0] operation_274_3898;
wire [7:0] operation_274_3897;
wire [7:0] operation_274_3896;
wire [7:0] operation_274_3895;
wire [7:0] operation_274_5467;
wire [7:0] operation_274_5466;
wire [7:0] operation_274_5465;
wire [7:0] operation_274_5444;
reg signed [31:0] operation_274_3927;
reg signed [31:0] operation_274_3926;
reg signed [31:0] operation_274_3925;
reg signed [31:0] operation_274_3924;
reg signed [31:0] operation_274_3923;
reg signed [31:0] operation_274_3922;
reg signed [31:0] operation_274_3921;
reg signed [31:0] operation_274_3920;
reg signed [31:0] operation_274_3919;
reg signed [31:0] operation_274_3918;
reg signed [31:0] operation_274_3917;
reg signed [31:0] operation_274_3916;
reg signed [31:0] operation_274_3915;
reg signed [31:0] operation_274_3914;
reg signed [31:0] operation_274_3913;
reg signed [31:0] operation_274_3912;
reg signed [31:0] operation_274_5488;
reg signed [31:0] operation_274_5487;
reg signed [31:0] operation_274_5486;
reg signed [31:0] operation_274_5469;
wire signed [31:0] operation_274_3945;
wire signed [31:0] operation_274_3944;
wire signed [31:0] operation_274_3943;
wire signed [31:0] operation_274_3942;
wire signed [31:0] operation_274_3941;
wire signed [31:0] operation_274_3940;
wire signed [31:0] operation_274_3939;
wire signed [31:0] operation_274_3938;
wire signed [31:0] operation_274_3937;
wire signed [31:0] operation_274_3936;
wire signed [31:0] operation_274_3935;
wire signed [31:0] operation_274_3934;
wire signed [31:0] operation_274_3933;
wire signed [31:0] operation_274_3932;
wire signed [31:0] operation_274_3931;
wire signed [31:0] operation_274_3930;
wire signed [31:0] operation_274_5510;
wire signed [31:0] operation_274_5509;
wire signed [31:0] operation_274_5508;
wire signed [31:0] operation_274_5491;
wire [7:0] operation_274_3965;
wire [7:0] operation_274_3964;
wire [7:0] operation_274_3963;
wire [7:0] operation_274_3962;
wire [7:0] operation_274_3961;
wire [7:0] operation_274_3960;
wire [7:0] operation_274_3959;
wire [7:0] operation_274_3958;
wire [7:0] operation_274_3957;
wire [7:0] operation_274_3956;
wire [7:0] operation_274_3955;
wire [7:0] operation_274_3954;
wire [7:0] operation_274_3953;
wire [7:0] operation_274_3952;
wire [7:0] operation_274_3951;
wire [7:0] operation_274_3950;
wire signed [31:0] operation_274_4805;
wire signed [31:0] operation_274_4804;
wire signed [31:0] operation_274_4786;
wire signed [31:0] operation_274_4735;
reg [7:0] operation_274_5538_latch;
wire [7:0] operation_274_5538;
reg [7:0] operation_274_5537_latch;
wire [7:0] operation_274_5537;
reg [7:0] operation_274_5520_latch;
wire [7:0] operation_274_5520;
reg [7:0] operation_274_5519_latch;
wire [7:0] operation_274_5519;
reg signed [31:0] operation_274_3985;
reg signed [31:0] operation_274_3984;
reg signed [31:0] operation_274_3983;
reg signed [31:0] operation_274_3982;
reg signed [31:0] operation_274_3981;
reg signed [31:0] operation_274_3980;
reg signed [31:0] operation_274_3979;
reg signed [31:0] operation_274_3978;
reg signed [31:0] operation_274_3977;
reg signed [31:0] operation_274_3976;
reg signed [31:0] operation_274_3975;
reg signed [31:0] operation_274_3974;
reg signed [31:0] operation_274_3973;
reg signed [31:0] operation_274_3972;
reg signed [31:0] operation_274_3971;
reg signed [31:0] operation_274_3970;
wire [7:0] operation_274_4825;
wire [7:0] operation_274_4824;
wire [7:0] operation_274_4806;
wire [7:0] operation_274_4752;
wire signed [31:0] operation_274_4005;
wire signed [31:0] operation_274_4004;
wire signed [31:0] operation_274_4003;
wire signed [31:0] operation_274_4002;
wire signed [31:0] operation_274_4001;
wire signed [31:0] operation_274_4000;
wire signed [31:0] operation_274_3999;
wire signed [31:0] operation_274_3998;
wire signed [31:0] operation_274_3997;
wire signed [31:0] operation_274_3996;
wire signed [31:0] operation_274_3995;
wire signed [31:0] operation_274_3994;
wire signed [31:0] operation_274_3993;
wire signed [31:0] operation_274_3992;
wire signed [31:0] operation_274_3991;
wire signed [31:0] operation_274_3990;
reg signed [31:0] operation_274_4845;
reg signed [31:0] operation_274_4844;
reg signed [31:0] operation_274_4826;
reg signed [31:0] operation_274_4769;
wire [7:0] operation_274_4025;
wire [7:0] operation_274_4024;
wire [7:0] operation_274_4023;
wire [7:0] operation_274_4022;
wire [7:0] operation_274_4021;
wire [7:0] operation_274_4020;
wire [7:0] operation_274_4019;
wire [7:0] operation_274_4018;
wire [7:0] operation_274_4017;
wire [7:0] operation_274_4016;
wire [7:0] operation_274_4015;
wire [7:0] operation_274_4014;
wire [7:0] operation_274_4013;
wire [7:0] operation_274_4012;
wire [7:0] operation_274_4011;
wire [7:0] operation_274_4010;
wire signed [31:0] operation_274_4865;
wire signed [31:0] operation_274_4864;
wire signed [31:0] operation_274_4846;
wire signed [31:0] operation_274_4787;
reg signed [31:0] operation_274_4045;
reg signed [31:0] operation_274_4044;
reg signed [31:0] operation_274_4043;
reg signed [31:0] operation_274_4042;
reg signed [31:0] operation_274_4041;
reg signed [31:0] operation_274_4040;
reg signed [31:0] operation_274_4039;
reg signed [31:0] operation_274_4038;
reg signed [31:0] operation_274_4037;
reg signed [31:0] operation_274_4036;
reg signed [31:0] operation_274_4035;
reg signed [31:0] operation_274_4034;
reg signed [31:0] operation_274_4033;
reg signed [31:0] operation_274_4032;
reg signed [31:0] operation_274_4031;
reg signed [31:0] operation_274_4030;
wire [7:0] operation_274_4885;
wire [7:0] operation_274_4884;
wire [7:0] operation_274_4866;
wire [7:0] operation_274_4807;
reg signed [31:0] operation_274_4065;
reg signed [31:0] operation_274_4064;
reg signed [31:0] operation_274_4063;
reg signed [31:0] operation_274_4062;
reg signed [31:0] operation_274_4061;
reg signed [31:0] operation_274_4060;
reg signed [31:0] operation_274_4059;
reg signed [31:0] operation_274_4058;
reg signed [31:0] operation_274_4057;
reg signed [31:0] operation_274_4056;
reg signed [31:0] operation_274_4055;
reg signed [31:0] operation_274_4054;
reg signed [31:0] operation_274_4053;
reg signed [31:0] operation_274_4052;
reg signed [31:0] operation_274_4051;
reg signed [31:0] operation_274_4050;
reg signed [31:0] operation_274_4905;
reg signed [31:0] operation_274_4904;
reg signed [31:0] operation_274_4886;
reg signed [31:0] operation_274_4827;
reg signed [31:0] operation_274_4089;
reg signed [31:0] operation_274_4088;
reg signed [31:0] operation_274_4087;
reg signed [31:0] operation_274_4086;
reg signed [31:0] operation_274_4085;
reg signed [31:0] operation_274_4084;
reg signed [31:0] operation_274_4083;
reg signed [31:0] operation_274_4082;
reg signed [31:0] operation_274_4081;
reg signed [31:0] operation_274_4080;
reg signed [31:0] operation_274_4079;
reg signed [31:0] operation_274_4078;
reg signed [31:0] operation_274_4077;
reg signed [31:0] operation_274_4076;
reg signed [31:0] operation_274_4075;
reg signed [31:0] operation_274_4074;
wire signed [31:0] operation_274_4073;
wire signed [31:0] operation_274_4072;
wire signed [31:0] operation_274_4071;
wire signed [31:0] operation_274_4070;
wire signed [31:0] operation_274_4925;
wire signed [31:0] operation_274_4924;
wire signed [31:0] operation_274_4906;
wire signed [31:0] operation_274_4847;
wire [7:0] operation_274_4129;
wire [7:0] operation_274_4128;
reg signed [31:0] operation_274_4127;
reg signed [31:0] operation_274_4126;
reg signed [31:0] operation_274_4125;
reg signed [31:0] operation_274_4124;
reg signed [31:0] operation_274_4123;
reg signed [31:0] operation_274_4122;
reg signed [31:0] operation_274_4121;
reg signed [31:0] operation_274_4120;
reg signed [31:0] operation_274_4119;
reg signed [31:0] operation_274_4118;
reg signed [31:0] operation_274_4117;
reg signed [31:0] operation_274_4116;
reg signed [31:0] operation_274_4115;
reg signed [31:0] operation_274_4114;
reg signed [31:0] operation_274_4113;
reg signed [31:0] operation_274_4112;
reg signed [31:0] operation_274_4111;
reg signed [31:0] operation_274_4110;
reg signed [31:0] operation_274_4109;
reg signed [31:0] operation_274_4108;
reg signed [31:0] operation_274_4107;
reg signed [31:0] operation_274_4106;
reg signed [31:0] operation_274_4105;
reg signed [31:0] operation_274_4104;
reg signed [31:0] operation_274_4103;
reg signed [31:0] operation_274_4102;
reg signed [31:0] operation_274_4101;
reg signed [31:0] operation_274_4100;
reg signed [31:0] operation_274_4099;
reg signed [31:0] operation_274_4098;
reg signed [31:0] operation_274_4097;
reg signed [31:0] operation_274_4096;
wire [7:0] operation_274_4095;
wire [7:0] operation_274_4094;
wire [7:0] operation_274_4949;
wire [7:0] operation_274_4948;
wire [7:0] operation_274_4926;
wire [7:0] operation_274_4867;
reg signed [31:0] operation_274_4153;
reg signed [31:0] operation_274_4152;
wire signed [31:0] operation_274_4151;
wire signed [31:0] operation_274_4150;
wire signed [31:0] operation_274_4149;
wire signed [31:0] operation_274_4148;
wire signed [31:0] operation_274_4147;
wire signed [31:0] operation_274_4146;
wire signed [31:0] operation_274_4145;
wire signed [31:0] operation_274_4144;
wire signed [31:0] operation_274_4143;
wire signed [31:0] operation_274_4142;
wire signed [31:0] operation_274_4141;
wire signed [31:0] operation_274_4140;
wire signed [31:0] operation_274_4139;
wire signed [31:0] operation_274_4138;
wire signed [31:0] operation_274_4137;
wire signed [31:0] operation_274_4136;
reg signed [31:0] operation_274_4135;
reg signed [31:0] operation_274_4134;
reg signed [31:0] operation_274_4989;
reg signed [31:0] operation_274_4988;
reg signed [31:0] operation_274_4950;
reg signed [31:0] operation_274_4887;
reg signed [31:0] operation_274_4177;
reg signed [31:0] operation_274_4176;
wire [7:0] operation_274_4175;
wire [7:0] operation_274_4174;
wire [7:0] operation_274_4173;
wire [7:0] operation_274_4172;
wire [7:0] operation_274_4171;
wire [7:0] operation_274_4170;
wire [7:0] operation_274_4169;
wire [7:0] operation_274_4168;
wire [7:0] operation_274_4167;
wire [7:0] operation_274_4166;
wire [7:0] operation_274_4165;
wire [7:0] operation_274_4164;
wire [7:0] operation_274_4163;
wire [7:0] operation_274_4162;
wire [7:0] operation_274_4161;
wire [7:0] operation_274_4160;
reg signed [31:0] operation_274_4159;
reg signed [31:0] operation_274_4158;
wire signed [31:0] operation_274_5013;
wire signed [31:0] operation_274_5012;
wire signed [31:0] operation_274_4990;
wire signed [31:0] operation_274_4907;
reg signed [31:0] operation_274_4198;
reg signed [31:0] operation_274_4197;
reg signed [31:0] operation_274_4196;
reg signed [31:0] operation_274_4195;
reg signed [31:0] operation_274_4194;
reg signed [31:0] operation_274_4193;
reg signed [31:0] operation_274_4192;
reg signed [31:0] operation_274_4191;
reg signed [31:0] operation_274_4190;
reg signed [31:0] operation_274_4189;
reg signed [31:0] operation_274_4188;
reg signed [31:0] operation_274_4187;
reg signed [31:0] operation_274_4186;
reg signed [31:0] operation_274_4185;
reg signed [31:0] operation_274_4184;
reg signed [31:0] operation_274_4183;
wire [7:0] operation_274_5038;
wire [7:0] operation_274_5037;
wire [7:0] operation_274_5015;
wire [7:0] operation_274_4927;
wire signed [31:0] operation_274_4220;
wire signed [31:0] operation_274_4219;
wire signed [31:0] operation_274_4218;
wire signed [31:0] operation_274_4217;
wire signed [31:0] operation_274_4216;
wire signed [31:0] operation_274_4215;
wire signed [31:0] operation_274_4214;
wire signed [31:0] operation_274_4213;
wire signed [31:0] operation_274_4212;
wire signed [31:0] operation_274_4211;
wire signed [31:0] operation_274_4210;
wire signed [31:0] operation_274_4209;
wire signed [31:0] operation_274_4208;
wire signed [31:0] operation_274_4207;
wire signed [31:0] operation_274_4206;
wire signed [31:0] operation_274_4205;
reg signed [31:0] operation_274_5059;
reg signed [31:0] operation_274_5058;
reg signed [31:0] operation_274_5040;
reg signed [31:0] operation_274_4951;
reg [7:0] operation_274_4249_latch;
wire [7:0] operation_274_4249;
reg [7:0] operation_274_4248_latch;
wire [7:0] operation_274_4248;
reg [7:0] operation_274_4247_latch;
wire [7:0] operation_274_4247;
reg [7:0] operation_274_4246_latch;
wire [7:0] operation_274_4246;
reg [7:0] operation_274_4245_latch;
wire [7:0] operation_274_4245;
reg [7:0] operation_274_4244_latch;
wire [7:0] operation_274_4244;
reg [7:0] operation_274_4243_latch;
wire [7:0] operation_274_4243;
reg [7:0] operation_274_4242_latch;
wire [7:0] operation_274_4242;
reg [7:0] operation_274_4241_latch;
wire [7:0] operation_274_4241;
reg [7:0] operation_274_4240_latch;
wire [7:0] operation_274_4240;
reg [7:0] operation_274_4239_latch;
wire [7:0] operation_274_4239;
reg [7:0] operation_274_4238_latch;
wire [7:0] operation_274_4238;
reg [7:0] operation_274_4237_latch;
wire [7:0] operation_274_4237;
reg [7:0] operation_274_4236_latch;
wire [7:0] operation_274_4236;
reg [7:0] operation_274_4235_latch;
wire [7:0] operation_274_4235;
reg [7:0] operation_274_4234_latch;
wire [7:0] operation_274_4234;
wire signed [31:0] operation_274_5081;
wire signed [31:0] operation_274_5080;
wire signed [31:0] operation_274_5062;
wire signed [31:0] operation_274_4991;
wire [7:0] operation_274_3430;
wire [7:0] operation_274_3429;
wire [7:0] operation_274_3428;
wire [7:0] operation_274_3427;
wire [7:0] operation_274_3426;
wire [7:0] operation_274_3425;
wire [7:0] operation_274_3424;
wire [7:0] operation_274_3423;
wire [7:0] operation_274_3422;
wire [7:0] operation_274_3421;
wire [7:0] operation_274_3420;
wire [7:0] operation_274_3419;
wire [7:0] operation_274_3418;
wire [7:0] operation_274_3417;
wire [7:0] operation_274_3416;
wire [7:0] operation_274_3415;
wire signed [31:0] operation_274_4376;
wire signed [31:0] operation_274_4357;
wire signed [31:0] operation_274_4306;
reg [7:0] operation_274_5109_latch;
wire [7:0] operation_274_5109;
reg [7:0] operation_274_5091_latch;
wire [7:0] operation_274_5091;
reg [7:0] operation_274_5090_latch;
wire [7:0] operation_274_5090;
wire [7:0] operation_274_5036;
reg signed [31:0] operation_274_3446;
reg signed [31:0] operation_274_3445;
reg signed [31:0] operation_274_3444;
reg signed [31:0] operation_274_3443;
reg signed [31:0] operation_274_3442;
reg signed [31:0] operation_274_3441;
reg signed [31:0] operation_274_3440;
reg signed [31:0] operation_274_3439;
reg signed [31:0] operation_274_3438;
reg signed [31:0] operation_274_3437;
reg signed [31:0] operation_274_3436;
reg signed [31:0] operation_274_3435;
reg signed [31:0] operation_274_3434;
reg signed [31:0] operation_274_3433;
reg signed [31:0] operation_274_3432;
reg signed [31:0] operation_274_3431;
wire [7:0] operation_274_4396;
wire [7:0] operation_274_4377;
wire [7:0] operation_274_4323;
reg signed [31:0] operation_274_5057;
wire signed [31:0] operation_274_3464;
wire signed [31:0] operation_274_3463;
wire signed [31:0] operation_274_3462;
wire signed [31:0] operation_274_3461;
wire signed [31:0] operation_274_3460;
wire signed [31:0] operation_274_3459;
wire signed [31:0] operation_274_3458;
wire signed [31:0] operation_274_3457;
wire signed [31:0] operation_274_3455;
wire signed [31:0] operation_274_3454;
wire signed [31:0] operation_274_3453;
wire signed [31:0] operation_274_3452;
wire signed [31:0] operation_274_3451;
wire signed [31:0] operation_274_3450;
wire signed [31:0] operation_274_3449;
wire signed [31:0] operation_274_3447;
reg signed [31:0] operation_274_4416;
reg signed [31:0] operation_274_4397;
reg signed [31:0] operation_274_4340;
wire signed [31:0] operation_274_5079;
wire [7:0] operation_274_3481;
wire [7:0] operation_274_3480;
wire [7:0] operation_274_3479;
wire [7:0] operation_274_3478;
wire [7:0] operation_274_3477;
wire [7:0] operation_274_3476;
wire [7:0] operation_274_3475;
wire [7:0] operation_274_3474;
wire [7:0] operation_274_3473;
wire [7:0] operation_274_3472;
wire [7:0] operation_274_3471;
wire [7:0] operation_274_3470;
wire [7:0] operation_274_3469;
wire [7:0] operation_274_3468;
wire [7:0] operation_274_3467;
wire [7:0] operation_274_3466;
wire signed [31:0] operation_274_4436;
wire signed [31:0] operation_274_4417;
wire signed [31:0] operation_274_4375;
wire signed [31:0] operation_274_4358;
reg [7:0] operation_274_5108_latch;
wire [7:0] operation_274_5108;
reg signed [31:0] operation_274_3498;
reg signed [31:0] operation_274_3497;
reg signed [31:0] operation_274_3496;
reg signed [31:0] operation_274_3495;
reg signed [31:0] operation_274_3494;
reg signed [31:0] operation_274_3493;
reg signed [31:0] operation_274_3492;
reg signed [31:0] operation_274_3491;
reg signed [31:0] operation_274_3490;
reg signed [31:0] operation_274_3489;
reg signed [31:0] operation_274_3488;
reg signed [31:0] operation_274_3487;
reg signed [31:0] operation_274_3486;
reg signed [31:0] operation_274_3485;
reg signed [31:0] operation_274_3484;
reg signed [31:0] operation_274_3483;
wire [7:0] operation_274_4456;
wire [7:0] operation_274_4437;
wire [7:0] operation_274_4395;
wire [7:0] operation_274_4378;
wire signed [31:0] operation_274_3516;
wire signed [31:0] operation_274_3515;
wire signed [31:0] operation_274_3514;
wire signed [31:0] operation_274_3513;
wire signed [31:0] operation_274_3512;
wire signed [31:0] operation_274_3511;
wire signed [31:0] operation_274_3510;
wire signed [31:0] operation_274_3509;
wire signed [31:0] operation_274_3508;
wire signed [31:0] operation_274_3507;
wire signed [31:0] operation_274_3506;
wire signed [31:0] operation_274_3505;
wire signed [31:0] operation_274_3504;
wire signed [31:0] operation_274_3503;
wire signed [31:0] operation_274_3502;
wire signed [31:0] operation_274_3501;
reg signed [31:0] operation_274_4476;
reg signed [31:0] operation_274_4457;
reg signed [31:0] operation_274_4415;
reg signed [31:0] operation_274_4398;
wire [7:0] operation_274_3536;
wire [7:0] operation_274_3535;
wire [7:0] operation_274_3534;
wire [7:0] operation_274_3533;
wire [7:0] operation_274_3532;
wire [7:0] operation_274_3531;
wire [7:0] operation_274_3530;
wire [7:0] operation_274_3529;
wire [7:0] operation_274_3528;
wire [7:0] operation_274_3527;
wire [7:0] operation_274_3526;
wire [7:0] operation_274_3525;
wire [7:0] operation_274_3524;
wire [7:0] operation_274_3523;
wire [7:0] operation_274_3522;
wire [7:0] operation_274_3521;
wire signed [31:0] operation_274_4496;
wire signed [31:0] operation_274_4477;
wire signed [31:0] operation_274_4435;
wire signed [31:0] operation_274_4418;
reg signed [31:0] operation_274_3556;
reg signed [31:0] operation_274_3555;
reg signed [31:0] operation_274_3554;
reg signed [31:0] operation_274_3553;
reg signed [31:0] operation_274_3552;
reg signed [31:0] operation_274_3551;
reg signed [31:0] operation_274_3550;
reg signed [31:0] operation_274_3549;
reg signed [31:0] operation_274_3548;
reg signed [31:0] operation_274_3547;
reg signed [31:0] operation_274_3546;
reg signed [31:0] operation_274_3545;
reg signed [31:0] operation_274_3544;
reg signed [31:0] operation_274_3543;
reg signed [31:0] operation_274_3542;
reg signed [31:0] operation_274_3541;
wire [7:0] operation_274_4520;
wire [7:0] operation_274_4497;
wire [7:0] operation_274_4455;
wire [7:0] operation_274_4438;
wire signed [31:0] operation_274_3576;
wire signed [31:0] operation_274_3575;
wire signed [31:0] operation_274_3574;
wire signed [31:0] operation_274_3573;
wire signed [31:0] operation_274_3572;
wire signed [31:0] operation_274_3571;
wire signed [31:0] operation_274_3570;
wire signed [31:0] operation_274_3569;
wire signed [31:0] operation_274_3568;
wire signed [31:0] operation_274_3567;
wire signed [31:0] operation_274_3566;
wire signed [31:0] operation_274_3565;
wire signed [31:0] operation_274_3564;
wire signed [31:0] operation_274_3563;
wire signed [31:0] operation_274_3562;
wire signed [31:0] operation_274_3561;
reg signed [31:0] operation_274_4560;
reg signed [31:0] operation_274_4521;
reg signed [31:0] operation_274_4475;
reg signed [31:0] operation_274_4458;
wire [7:0] operation_274_3596;
wire [7:0] operation_274_3595;
wire [7:0] operation_274_3594;
wire [7:0] operation_274_3593;
wire [7:0] operation_274_3592;
wire [7:0] operation_274_3591;
wire [7:0] operation_274_3590;
wire [7:0] operation_274_3589;
wire [7:0] operation_274_3588;
wire [7:0] operation_274_3587;
wire [7:0] operation_274_3586;
wire [7:0] operation_274_3585;
wire [7:0] operation_274_3584;
wire [7:0] operation_274_3583;
wire [7:0] operation_274_3582;
wire [7:0] operation_274_3581;
wire signed [31:0] operation_274_4584;
wire signed [31:0] operation_274_4561;
wire signed [31:0] operation_274_4495;
wire signed [31:0] operation_274_4478;
reg signed [31:0] operation_274_3616;
reg signed [31:0] operation_274_3615;
reg signed [31:0] operation_274_3614;
reg signed [31:0] operation_274_3613;
reg signed [31:0] operation_274_3612;
reg signed [31:0] operation_274_3611;
reg signed [31:0] operation_274_3610;
reg signed [31:0] operation_274_3609;
reg signed [31:0] operation_274_3608;
reg signed [31:0] operation_274_3607;
reg signed [31:0] operation_274_3606;
reg signed [31:0] operation_274_3605;
reg signed [31:0] operation_274_3604;
reg signed [31:0] operation_274_3603;
reg signed [31:0] operation_274_3602;
reg signed [31:0] operation_274_3601;
wire [7:0] operation_274_4609;
wire [7:0] operation_274_4586;
wire [7:0] operation_274_4519;
wire [7:0] operation_274_4498;
reg signed [31:0] operation_274_3636;
reg signed [31:0] operation_274_3635;
reg signed [31:0] operation_274_3634;
reg signed [31:0] operation_274_3633;
reg signed [31:0] operation_274_3632;
reg signed [31:0] operation_274_3631;
reg signed [31:0] operation_274_3630;
reg signed [31:0] operation_274_3629;
reg signed [31:0] operation_274_3628;
reg signed [31:0] operation_274_3627;
reg signed [31:0] operation_274_3626;
reg signed [31:0] operation_274_3625;
reg signed [31:0] operation_274_3624;
reg signed [31:0] operation_274_3623;
reg signed [31:0] operation_274_3622;
reg signed [31:0] operation_274_3621;
reg signed [31:0] operation_274_4630;
reg signed [31:0] operation_274_4611;
reg signed [31:0] operation_274_4559;
reg signed [31:0] operation_274_4522;
reg signed [31:0] operation_274_3660;
reg signed [31:0] operation_274_3659;
reg signed [31:0] operation_274_3658;
reg signed [31:0] operation_274_3657;
reg signed [31:0] operation_274_3656;
reg signed [31:0] operation_274_3655;
reg signed [31:0] operation_274_3654;
reg signed [31:0] operation_274_3653;
reg signed [31:0] operation_274_3652;
reg signed [31:0] operation_274_3651;
reg signed [31:0] operation_274_3650;
reg signed [31:0] operation_274_3649;
reg signed [31:0] operation_274_3648;
reg signed [31:0] operation_274_3647;
reg signed [31:0] operation_274_3646;
reg signed [31:0] operation_274_3645;
wire signed [31:0] operation_274_3644;
wire signed [31:0] operation_274_3643;
wire signed [31:0] operation_274_3642;
wire signed [31:0] operation_274_3641;
wire signed [31:0] operation_274_4652;
wire signed [31:0] operation_274_4633;
wire signed [31:0] operation_274_4583;
wire signed [31:0] operation_274_4562;
wire [7:0] operation_274_3700;
wire [7:0] operation_274_3699;
reg signed [31:0] operation_274_3698;
reg signed [31:0] operation_274_3697;
reg signed [31:0] operation_274_3696;
reg signed [31:0] operation_274_3695;
reg signed [31:0] operation_274_3694;
reg signed [31:0] operation_274_3693;
reg signed [31:0] operation_274_3692;
reg signed [31:0] operation_274_3691;
reg signed [31:0] operation_274_3690;
reg signed [31:0] operation_274_3689;
reg signed [31:0] operation_274_3688;
reg signed [31:0] operation_274_3687;
reg signed [31:0] operation_274_3686;
reg signed [31:0] operation_274_3685;
reg signed [31:0] operation_274_3684;
reg signed [31:0] operation_274_3683;
reg signed [31:0] operation_274_3682;
reg signed [31:0] operation_274_3681;
reg signed [31:0] operation_274_3680;
reg signed [31:0] operation_274_3679;
reg signed [31:0] operation_274_3678;
reg signed [31:0] operation_274_3677;
reg signed [31:0] operation_274_3676;
reg signed [31:0] operation_274_3675;
reg signed [31:0] operation_274_3674;
reg signed [31:0] operation_274_3673;
reg signed [31:0] operation_274_3672;
reg signed [31:0] operation_274_3671;
reg signed [31:0] operation_274_3670;
reg signed [31:0] operation_274_3669;
reg signed [31:0] operation_274_3668;
reg signed [31:0] operation_274_3667;
wire [7:0] operation_274_3666;
wire [7:0] operation_274_3665;
wire signed [31:0] operation_274_3947;
wire signed [31:0] operation_274_3877;
reg [7:0] operation_274_4680_latch;
wire [7:0] operation_274_4680;
reg [7:0] operation_274_4661_latch;
wire [7:0] operation_274_4661;
wire [7:0] operation_274_4608;
wire [7:0] operation_274_4607;
reg signed [31:0] operation_274_3724;
reg signed [31:0] operation_274_3723;
wire signed [31:0] operation_274_3722;
wire signed [31:0] operation_274_3721;
wire signed [31:0] operation_274_3720;
wire signed [31:0] operation_274_3719;
wire signed [31:0] operation_274_3718;
wire signed [31:0] operation_274_3717;
wire signed [31:0] operation_274_3716;
wire signed [31:0] operation_274_3715;
wire signed [31:0] operation_274_3714;
wire signed [31:0] operation_274_3713;
wire signed [31:0] operation_274_3712;
wire signed [31:0] operation_274_3711;
wire signed [31:0] operation_274_3710;
wire signed [31:0] operation_274_3709;
wire signed [31:0] operation_274_3708;
wire signed [31:0] operation_274_3707;
reg signed [31:0] operation_274_3706;
reg signed [31:0] operation_274_3705;
wire [7:0] operation_274_3967;
wire [7:0] operation_274_3894;
reg signed [31:0] operation_274_4629;
reg signed [31:0] operation_274_4628;
reg signed [31:0] operation_274_3748;
reg signed [31:0] operation_274_3747;
wire [7:0] operation_274_3746;
wire [7:0] operation_274_3745;
wire [7:0] operation_274_3744;
wire [7:0] operation_274_3743;
wire [7:0] operation_274_3742;
wire [7:0] operation_274_3741;
wire [7:0] operation_274_3740;
wire [7:0] operation_274_3739;
wire [7:0] operation_274_3738;
wire [7:0] operation_274_3737;
wire [7:0] operation_274_3736;
wire [7:0] operation_274_3735;
wire [7:0] operation_274_3734;
wire [7:0] operation_274_3733;
wire [7:0] operation_274_3732;
wire [7:0] operation_274_3731;
reg signed [31:0] operation_274_3730;
reg signed [31:0] operation_274_3729;
reg signed [31:0] operation_274_3987;
reg signed [31:0] operation_274_3911;
wire signed [31:0] operation_274_4651;
wire signed [31:0] operation_274_4650;
reg signed [31:0] operation_274_3769;
reg signed [31:0] operation_274_3768;
reg signed [31:0] operation_274_3767;
reg signed [31:0] operation_274_3766;
reg signed [31:0] operation_274_3765;
reg signed [31:0] operation_274_3764;
reg signed [31:0] operation_274_3763;
reg signed [31:0] operation_274_3762;
reg signed [31:0] operation_274_3761;
reg signed [31:0] operation_274_3760;
reg signed [31:0] operation_274_3759;
reg signed [31:0] operation_274_3758;
reg signed [31:0] operation_274_3757;
reg signed [31:0] operation_274_3756;
reg signed [31:0] operation_274_3755;
reg signed [31:0] operation_274_3754;
wire signed [31:0] operation_274_4007;
wire signed [31:0] operation_274_3946;
wire signed [31:0] operation_274_3929;
wire signed [31:0] operation_274_3928;
reg [7:0] operation_274_4679_latch;
wire [7:0] operation_274_4679;
reg [7:0] operation_274_4662_latch;
wire [7:0] operation_274_4662;
wire signed [31:0] operation_274_3791;
wire signed [31:0] operation_274_3790;
wire signed [31:0] operation_274_3789;
wire signed [31:0] operation_274_3788;
wire signed [31:0] operation_274_3787;
wire signed [31:0] operation_274_3786;
wire signed [31:0] operation_274_3785;
wire signed [31:0] operation_274_3784;
wire signed [31:0] operation_274_3783;
wire signed [31:0] operation_274_3782;
wire signed [31:0] operation_274_3781;
wire signed [31:0] operation_274_3780;
wire signed [31:0] operation_274_3779;
wire signed [31:0] operation_274_3778;
wire signed [31:0] operation_274_3777;
wire signed [31:0] operation_274_3776;
wire [7:0] operation_274_4027;
wire [7:0] operation_274_3966;
wire [7:0] operation_274_3949;
wire [7:0] operation_274_3948;
reg [7:0] operation_274_3820_latch;
wire [7:0] operation_274_3820;
reg [7:0] operation_274_3819_latch;
wire [7:0] operation_274_3819;
reg [7:0] operation_274_3818_latch;
wire [7:0] operation_274_3818;
reg [7:0] operation_274_3817_latch;
wire [7:0] operation_274_3817;
reg [7:0] operation_274_3816_latch;
wire [7:0] operation_274_3816;
reg [7:0] operation_274_3815_latch;
wire [7:0] operation_274_3815;
reg [7:0] operation_274_3814_latch;
wire [7:0] operation_274_3814;
reg [7:0] operation_274_3813_latch;
wire [7:0] operation_274_3813;
reg [7:0] operation_274_3812_latch;
wire [7:0] operation_274_3812;
reg [7:0] operation_274_3811_latch;
wire [7:0] operation_274_3811;
reg [7:0] operation_274_3810_latch;
wire [7:0] operation_274_3810;
reg [7:0] operation_274_3809_latch;
wire [7:0] operation_274_3809;
reg [7:0] operation_274_3808_latch;
wire [7:0] operation_274_3808;
reg [7:0] operation_274_3807_latch;
wire [7:0] operation_274_3807;
reg [7:0] operation_274_3806_latch;
wire [7:0] operation_274_3806;
reg [7:0] operation_274_3805_latch;
wire [7:0] operation_274_3805;
reg signed [31:0] operation_274_4047;
reg signed [31:0] operation_274_3986;
reg signed [31:0] operation_274_3969;
reg signed [31:0] operation_274_3968;
wire [7:0] operation_274_3001;
wire [7:0] operation_274_3000;
wire [7:0] operation_274_2999;
wire [7:0] operation_274_2998;
wire [7:0] operation_274_2997;
wire [7:0] operation_274_2996;
wire [7:0] operation_274_2995;
wire [7:0] operation_274_2994;
wire [7:0] operation_274_2993;
wire [7:0] operation_274_2992;
wire [7:0] operation_274_2991;
wire [7:0] operation_274_2990;
wire [7:0] operation_274_2989;
wire [7:0] operation_274_2988;
wire [7:0] operation_274_2987;
wire [7:0] operation_274_2986;
wire signed [31:0] operation_274_4067;
wire signed [31:0] operation_274_4006;
wire signed [31:0] operation_274_3989;
wire signed [31:0] operation_274_3988;
reg signed [31:0] operation_274_3017;
reg signed [31:0] operation_274_3016;
reg signed [31:0] operation_274_3015;
reg signed [31:0] operation_274_3014;
reg signed [31:0] operation_274_3013;
reg signed [31:0] operation_274_3012;
reg signed [31:0] operation_274_3011;
reg signed [31:0] operation_274_3010;
reg signed [31:0] operation_274_3009;
reg signed [31:0] operation_274_3008;
reg signed [31:0] operation_274_3007;
reg signed [31:0] operation_274_3006;
reg signed [31:0] operation_274_3005;
reg signed [31:0] operation_274_3004;
reg signed [31:0] operation_274_3003;
reg signed [31:0] operation_274_3002;
wire [7:0] operation_274_4091;
wire [7:0] operation_274_4026;
wire [7:0] operation_274_4009;
wire [7:0] operation_274_4008;
wire signed [31:0] operation_274_3035;
wire signed [31:0] operation_274_3034;
wire signed [31:0] operation_274_3033;
wire signed [31:0] operation_274_3032;
wire signed [31:0] operation_274_3031;
wire signed [31:0] operation_274_3030;
wire signed [31:0] operation_274_3029;
wire signed [31:0] operation_274_3028;
wire signed [31:0] operation_274_3026;
wire signed [31:0] operation_274_3025;
wire signed [31:0] operation_274_3024;
wire signed [31:0] operation_274_3023;
wire signed [31:0] operation_274_3022;
wire signed [31:0] operation_274_3021;
wire signed [31:0] operation_274_3020;
wire signed [31:0] operation_274_3018;
reg signed [31:0] operation_274_4131;
reg signed [31:0] operation_274_4046;
reg signed [31:0] operation_274_4029;
reg signed [31:0] operation_274_4028;
wire [7:0] operation_274_3052;
wire [7:0] operation_274_3051;
wire [7:0] operation_274_3050;
wire [7:0] operation_274_3049;
wire [7:0] operation_274_3048;
wire [7:0] operation_274_3047;
wire [7:0] operation_274_3046;
wire [7:0] operation_274_3045;
wire [7:0] operation_274_3044;
wire [7:0] operation_274_3043;
wire [7:0] operation_274_3042;
wire [7:0] operation_274_3041;
wire [7:0] operation_274_3040;
wire [7:0] operation_274_3039;
wire [7:0] operation_274_3038;
wire [7:0] operation_274_3037;
wire signed [31:0] operation_274_4155;
wire signed [31:0] operation_274_4066;
wire signed [31:0] operation_274_4049;
wire signed [31:0] operation_274_4048;
reg signed [31:0] operation_274_3069;
reg signed [31:0] operation_274_3068;
reg signed [31:0] operation_274_3067;
reg signed [31:0] operation_274_3066;
reg signed [31:0] operation_274_3065;
reg signed [31:0] operation_274_3064;
reg signed [31:0] operation_274_3063;
reg signed [31:0] operation_274_3062;
reg signed [31:0] operation_274_3061;
reg signed [31:0] operation_274_3060;
reg signed [31:0] operation_274_3059;
reg signed [31:0] operation_274_3058;
reg signed [31:0] operation_274_3057;
reg signed [31:0] operation_274_3056;
reg signed [31:0] operation_274_3055;
reg signed [31:0] operation_274_3054;
wire [7:0] operation_274_4180;
wire [7:0] operation_274_4090;
wire [7:0] operation_274_4069;
wire [7:0] operation_274_4068;
wire signed [31:0] operation_274_3087;
wire signed [31:0] operation_274_3086;
wire signed [31:0] operation_274_3085;
wire signed [31:0] operation_274_3084;
wire signed [31:0] operation_274_3083;
wire signed [31:0] operation_274_3082;
wire signed [31:0] operation_274_3081;
wire signed [31:0] operation_274_3080;
wire signed [31:0] operation_274_3079;
wire signed [31:0] operation_274_3078;
wire signed [31:0] operation_274_3077;
wire signed [31:0] operation_274_3076;
wire signed [31:0] operation_274_3075;
wire signed [31:0] operation_274_3074;
wire signed [31:0] operation_274_3073;
wire signed [31:0] operation_274_3072;
reg signed [31:0] operation_274_4201;
reg signed [31:0] operation_274_4130;
reg signed [31:0] operation_274_4093;
reg signed [31:0] operation_274_4092;
wire [7:0] operation_274_3107;
wire [7:0] operation_274_3106;
wire [7:0] operation_274_3105;
wire [7:0] operation_274_3104;
wire [7:0] operation_274_3103;
wire [7:0] operation_274_3102;
wire [7:0] operation_274_3101;
wire [7:0] operation_274_3100;
wire [7:0] operation_274_3099;
wire [7:0] operation_274_3098;
wire [7:0] operation_274_3097;
wire [7:0] operation_274_3096;
wire [7:0] operation_274_3095;
wire [7:0] operation_274_3094;
wire [7:0] operation_274_3093;
wire [7:0] operation_274_3092;
wire signed [31:0] operation_274_4223;
wire signed [31:0] operation_274_4154;
wire signed [31:0] operation_274_4133;
wire signed [31:0] operation_274_4132;
reg signed [31:0] operation_274_3127;
reg signed [31:0] operation_274_3126;
reg signed [31:0] operation_274_3125;
reg signed [31:0] operation_274_3124;
reg signed [31:0] operation_274_3123;
reg signed [31:0] operation_274_3122;
reg signed [31:0] operation_274_3121;
reg signed [31:0] operation_274_3120;
reg signed [31:0] operation_274_3119;
reg signed [31:0] operation_274_3118;
reg signed [31:0] operation_274_3117;
reg signed [31:0] operation_274_3116;
reg signed [31:0] operation_274_3115;
reg signed [31:0] operation_274_3114;
reg signed [31:0] operation_274_3113;
reg signed [31:0] operation_274_3112;
wire signed [31:0] operation_274_3448;
reg [7:0] operation_274_4232_latch;
wire [7:0] operation_274_4232;
wire [7:0] operation_274_4179;
wire [7:0] operation_274_4178;
wire [7:0] operation_274_4157;
wire signed [31:0] operation_274_3147;
wire signed [31:0] operation_274_3146;
wire signed [31:0] operation_274_3145;
wire signed [31:0] operation_274_3144;
wire signed [31:0] operation_274_3143;
wire signed [31:0] operation_274_3142;
wire signed [31:0] operation_274_3141;
wire signed [31:0] operation_274_3140;
wire signed [31:0] operation_274_3139;
wire signed [31:0] operation_274_3138;
wire signed [31:0] operation_274_3137;
wire signed [31:0] operation_274_3136;
wire signed [31:0] operation_274_3135;
wire signed [31:0] operation_274_3134;
wire signed [31:0] operation_274_3133;
wire signed [31:0] operation_274_3132;
wire [7:0] operation_274_3465;
reg signed [31:0] operation_274_4200;
reg signed [31:0] operation_274_4199;
reg signed [31:0] operation_274_4182;
wire [7:0] operation_274_3167;
wire [7:0] operation_274_3166;
wire [7:0] operation_274_3165;
wire [7:0] operation_274_3164;
wire [7:0] operation_274_3163;
wire [7:0] operation_274_3162;
wire [7:0] operation_274_3161;
wire [7:0] operation_274_3160;
wire [7:0] operation_274_3159;
wire [7:0] operation_274_3158;
wire [7:0] operation_274_3157;
wire [7:0] operation_274_3156;
wire [7:0] operation_274_3155;
wire [7:0] operation_274_3154;
wire [7:0] operation_274_3153;
wire [7:0] operation_274_3152;
reg signed [31:0] operation_274_3482;
wire signed [31:0] operation_274_4222;
wire signed [31:0] operation_274_4221;
wire signed [31:0] operation_274_4204;
reg signed [31:0] operation_274_3187;
reg signed [31:0] operation_274_3186;
reg signed [31:0] operation_274_3185;
reg signed [31:0] operation_274_3184;
reg signed [31:0] operation_274_3183;
reg signed [31:0] operation_274_3182;
reg signed [31:0] operation_274_3181;
reg signed [31:0] operation_274_3180;
reg signed [31:0] operation_274_3179;
reg signed [31:0] operation_274_3178;
reg signed [31:0] operation_274_3177;
reg signed [31:0] operation_274_3176;
reg signed [31:0] operation_274_3175;
reg signed [31:0] operation_274_3174;
reg signed [31:0] operation_274_3173;
reg signed [31:0] operation_274_3172;
wire signed [31:0] operation_274_3518;
wire signed [31:0] operation_274_3517;
wire signed [31:0] operation_274_3500;
wire signed [31:0] operation_274_3499;
reg [7:0] operation_274_4251_latch;
wire [7:0] operation_274_4251;
reg [7:0] operation_274_4250_latch;
wire [7:0] operation_274_4250;
reg [7:0] operation_274_4233_latch;
wire [7:0] operation_274_4233;
reg signed [31:0] operation_274_3207;
reg signed [31:0] operation_274_3206;
reg signed [31:0] operation_274_3205;
reg signed [31:0] operation_274_3204;
reg signed [31:0] operation_274_3203;
reg signed [31:0] operation_274_3202;
reg signed [31:0] operation_274_3201;
reg signed [31:0] operation_274_3200;
reg signed [31:0] operation_274_3199;
reg signed [31:0] operation_274_3198;
reg signed [31:0] operation_274_3197;
reg signed [31:0] operation_274_3196;
reg signed [31:0] operation_274_3195;
reg signed [31:0] operation_274_3194;
reg signed [31:0] operation_274_3193;
reg signed [31:0] operation_274_3192;
wire [7:0] operation_274_3538;
wire [7:0] operation_274_3537;
wire [7:0] operation_274_3520;
wire [7:0] operation_274_3519;
reg signed [31:0] operation_274_3231;
reg signed [31:0] operation_274_3230;
reg signed [31:0] operation_274_3229;
reg signed [31:0] operation_274_3228;
reg signed [31:0] operation_274_3227;
reg signed [31:0] operation_274_3226;
reg signed [31:0] operation_274_3225;
reg signed [31:0] operation_274_3224;
reg signed [31:0] operation_274_3223;
reg signed [31:0] operation_274_3222;
reg signed [31:0] operation_274_3221;
reg signed [31:0] operation_274_3220;
reg signed [31:0] operation_274_3219;
reg signed [31:0] operation_274_3218;
reg signed [31:0] operation_274_3217;
reg signed [31:0] operation_274_3216;
wire signed [31:0] operation_274_3215;
wire signed [31:0] operation_274_3214;
wire signed [31:0] operation_274_3213;
wire signed [31:0] operation_274_3212;
reg signed [31:0] operation_274_3558;
reg signed [31:0] operation_274_3557;
reg signed [31:0] operation_274_3540;
reg signed [31:0] operation_274_3539;
wire [7:0] operation_274_3271;
wire [7:0] operation_274_3270;
reg signed [31:0] operation_274_3269;
reg signed [31:0] operation_274_3268;
reg signed [31:0] operation_274_3267;
reg signed [31:0] operation_274_3266;
reg signed [31:0] operation_274_3265;
reg signed [31:0] operation_274_3264;
reg signed [31:0] operation_274_3263;
reg signed [31:0] operation_274_3262;
reg signed [31:0] operation_274_3261;
reg signed [31:0] operation_274_3260;
reg signed [31:0] operation_274_3259;
reg signed [31:0] operation_274_3258;
reg signed [31:0] operation_274_3257;
reg signed [31:0] operation_274_3256;
reg signed [31:0] operation_274_3255;
reg signed [31:0] operation_274_3254;
reg signed [31:0] operation_274_3253;
reg signed [31:0] operation_274_3252;
reg signed [31:0] operation_274_3251;
reg signed [31:0] operation_274_3250;
reg signed [31:0] operation_274_3249;
reg signed [31:0] operation_274_3248;
reg signed [31:0] operation_274_3247;
reg signed [31:0] operation_274_3246;
reg signed [31:0] operation_274_3245;
reg signed [31:0] operation_274_3244;
reg signed [31:0] operation_274_3243;
reg signed [31:0] operation_274_3242;
reg signed [31:0] operation_274_3241;
reg signed [31:0] operation_274_3240;
reg signed [31:0] operation_274_3239;
reg signed [31:0] operation_274_3238;
wire [7:0] operation_274_3237;
wire [7:0] operation_274_3236;
wire signed [31:0] operation_274_3578;
wire signed [31:0] operation_274_3577;
wire signed [31:0] operation_274_3560;
wire signed [31:0] operation_274_3559;
reg signed [31:0] operation_274_3295;
reg signed [31:0] operation_274_3294;
wire signed [31:0] operation_274_3293;
wire signed [31:0] operation_274_3292;
wire signed [31:0] operation_274_3291;
wire signed [31:0] operation_274_3290;
wire signed [31:0] operation_274_3289;
wire signed [31:0] operation_274_3288;
wire signed [31:0] operation_274_3287;
wire signed [31:0] operation_274_3286;
wire signed [31:0] operation_274_3285;
wire signed [31:0] operation_274_3284;
wire signed [31:0] operation_274_3283;
wire signed [31:0] operation_274_3282;
wire signed [31:0] operation_274_3281;
wire signed [31:0] operation_274_3280;
wire signed [31:0] operation_274_3279;
wire signed [31:0] operation_274_3278;
reg signed [31:0] operation_274_3277;
reg signed [31:0] operation_274_3276;
wire [7:0] operation_274_3598;
wire [7:0] operation_274_3597;
wire [7:0] operation_274_3580;
wire [7:0] operation_274_3579;
reg signed [31:0] operation_274_3319;
reg signed [31:0] operation_274_3318;
wire [7:0] operation_274_3317;
wire [7:0] operation_274_3316;
wire [7:0] operation_274_3315;
wire [7:0] operation_274_3314;
wire [7:0] operation_274_3313;
wire [7:0] operation_274_3312;
wire [7:0] operation_274_3311;
wire [7:0] operation_274_3310;
wire [7:0] operation_274_3309;
wire [7:0] operation_274_3308;
wire [7:0] operation_274_3307;
wire [7:0] operation_274_3306;
wire [7:0] operation_274_3305;
wire [7:0] operation_274_3304;
wire [7:0] operation_274_3303;
wire [7:0] operation_274_3302;
reg signed [31:0] operation_274_3301;
reg signed [31:0] operation_274_3300;
reg signed [31:0] operation_274_3618;
reg signed [31:0] operation_274_3617;
reg signed [31:0] operation_274_3600;
reg signed [31:0] operation_274_3599;
reg signed [31:0] operation_274_3340;
reg signed [31:0] operation_274_3339;
reg signed [31:0] operation_274_3338;
reg signed [31:0] operation_274_3337;
reg signed [31:0] operation_274_3336;
reg signed [31:0] operation_274_3335;
reg signed [31:0] operation_274_3334;
reg signed [31:0] operation_274_3333;
reg signed [31:0] operation_274_3332;
reg signed [31:0] operation_274_3331;
reg signed [31:0] operation_274_3330;
reg signed [31:0] operation_274_3329;
reg signed [31:0] operation_274_3328;
reg signed [31:0] operation_274_3327;
reg signed [31:0] operation_274_3326;
reg signed [31:0] operation_274_3325;
wire signed [31:0] operation_274_3638;
wire signed [31:0] operation_274_3637;
wire signed [31:0] operation_274_3620;
wire signed [31:0] operation_274_3619;
wire signed [31:0] operation_274_3362;
wire signed [31:0] operation_274_3361;
wire signed [31:0] operation_274_3360;
wire signed [31:0] operation_274_3359;
wire signed [31:0] operation_274_3358;
wire signed [31:0] operation_274_3357;
wire signed [31:0] operation_274_3356;
wire signed [31:0] operation_274_3355;
wire signed [31:0] operation_274_3354;
wire signed [31:0] operation_274_3353;
wire signed [31:0] operation_274_3352;
wire signed [31:0] operation_274_3351;
wire signed [31:0] operation_274_3350;
wire signed [31:0] operation_274_3349;
wire signed [31:0] operation_274_3348;
wire signed [31:0] operation_274_3347;
wire [7:0] operation_274_3662;
wire [7:0] operation_274_3661;
wire [7:0] operation_274_3640;
wire [7:0] operation_274_3639;
reg [7:0] operation_274_3391_latch;
wire [7:0] operation_274_3391;
reg [7:0] operation_274_3390_latch;
wire [7:0] operation_274_3390;
reg [7:0] operation_274_3389_latch;
wire [7:0] operation_274_3389;
reg [7:0] operation_274_3388_latch;
wire [7:0] operation_274_3388;
reg [7:0] operation_274_3387_latch;
wire [7:0] operation_274_3387;
reg [7:0] operation_274_3386_latch;
wire [7:0] operation_274_3386;
reg [7:0] operation_274_3385_latch;
wire [7:0] operation_274_3385;
reg [7:0] operation_274_3384_latch;
wire [7:0] operation_274_3384;
reg [7:0] operation_274_3383_latch;
wire [7:0] operation_274_3383;
reg [7:0] operation_274_3382_latch;
wire [7:0] operation_274_3382;
reg [7:0] operation_274_3381_latch;
wire [7:0] operation_274_3381;
reg [7:0] operation_274_3380_latch;
wire [7:0] operation_274_3380;
reg [7:0] operation_274_3379_latch;
wire [7:0] operation_274_3379;
reg [7:0] operation_274_3378_latch;
wire [7:0] operation_274_3378;
reg [7:0] operation_274_3377_latch;
wire [7:0] operation_274_3377;
reg [7:0] operation_274_3376_latch;
wire [7:0] operation_274_3376;
reg signed [31:0] operation_274_3702;
reg signed [31:0] operation_274_3701;
reg signed [31:0] operation_274_3664;
reg signed [31:0] operation_274_3663;
wire [7:0] operation_274_2572;
wire [7:0] operation_274_2571;
wire [7:0] operation_274_2570;
wire [7:0] operation_274_2569;
wire [7:0] operation_274_2568;
wire [7:0] operation_274_2567;
wire [7:0] operation_274_2566;
wire [7:0] operation_274_2565;
wire [7:0] operation_274_2564;
wire [7:0] operation_274_2563;
wire [7:0] operation_274_2562;
wire [7:0] operation_274_2561;
wire [7:0] operation_274_2560;
wire [7:0] operation_274_2559;
wire [7:0] operation_274_2558;
wire [7:0] operation_274_2557;
wire signed [31:0] operation_274_3726;
wire signed [31:0] operation_274_3725;
wire signed [31:0] operation_274_3704;
wire signed [31:0] operation_274_3703;
reg signed [31:0] operation_274_2588;
reg signed [31:0] operation_274_2587;
reg signed [31:0] operation_274_2586;
reg signed [31:0] operation_274_2585;
reg signed [31:0] operation_274_2584;
reg signed [31:0] operation_274_2583;
reg signed [31:0] operation_274_2582;
reg signed [31:0] operation_274_2581;
reg signed [31:0] operation_274_2580;
reg signed [31:0] operation_274_2579;
reg signed [31:0] operation_274_2578;
reg signed [31:0] operation_274_2577;
reg signed [31:0] operation_274_2576;
reg signed [31:0] operation_274_2575;
reg signed [31:0] operation_274_2574;
reg signed [31:0] operation_274_2573;
wire [7:0] operation_274_3751;
wire [7:0] operation_274_3750;
wire [7:0] operation_274_3749;
wire [7:0] operation_274_3728;
wire signed [31:0] operation_274_2606;
wire signed [31:0] operation_274_2605;
wire signed [31:0] operation_274_2604;
wire signed [31:0] operation_274_2603;
wire signed [31:0] operation_274_2602;
wire signed [31:0] operation_274_2601;
wire signed [31:0] operation_274_2600;
wire signed [31:0] operation_274_2599;
wire signed [31:0] operation_274_2597;
wire signed [31:0] operation_274_2596;
wire signed [31:0] operation_274_2595;
wire signed [31:0] operation_274_2594;
wire signed [31:0] operation_274_2593;
wire signed [31:0] operation_274_2592;
wire signed [31:0] operation_274_2591;
wire signed [31:0] operation_274_2589;
reg signed [31:0] operation_274_3772;
reg signed [31:0] operation_274_3771;
reg signed [31:0] operation_274_3770;
reg signed [31:0] operation_274_3753;
wire [7:0] operation_274_2623;
wire [7:0] operation_274_2622;
wire [7:0] operation_274_2621;
wire [7:0] operation_274_2620;
wire [7:0] operation_274_2619;
wire [7:0] operation_274_2618;
wire [7:0] operation_274_2617;
wire [7:0] operation_274_2616;
wire [7:0] operation_274_2615;
wire [7:0] operation_274_2614;
wire [7:0] operation_274_2613;
wire [7:0] operation_274_2612;
wire [7:0] operation_274_2611;
wire [7:0] operation_274_2610;
wire [7:0] operation_274_2609;
wire [7:0] operation_274_2608;
wire signed [31:0] operation_274_3794;
wire signed [31:0] operation_274_3793;
wire signed [31:0] operation_274_3792;
wire signed [31:0] operation_274_3775;
reg signed [31:0] operation_274_2640;
reg signed [31:0] operation_274_2639;
reg signed [31:0] operation_274_2638;
reg signed [31:0] operation_274_2637;
reg signed [31:0] operation_274_2636;
reg signed [31:0] operation_274_2635;
reg signed [31:0] operation_274_2634;
reg signed [31:0] operation_274_2633;
reg signed [31:0] operation_274_2632;
reg signed [31:0] operation_274_2631;
reg signed [31:0] operation_274_2630;
reg signed [31:0] operation_274_2629;
reg signed [31:0] operation_274_2628;
reg signed [31:0] operation_274_2627;
reg signed [31:0] operation_274_2626;
reg signed [31:0] operation_274_2625;
wire signed [31:0] operation_274_3089;
wire signed [31:0] operation_274_3088;
wire signed [31:0] operation_274_3070;
wire signed [31:0] operation_274_3019;
reg [7:0] operation_274_3822_latch;
wire [7:0] operation_274_3822;
reg [7:0] operation_274_3821_latch;
wire [7:0] operation_274_3821;
reg [7:0] operation_274_3804_latch;
wire [7:0] operation_274_3804;
reg [7:0] operation_274_3803_latch;
wire [7:0] operation_274_3803;
wire signed [31:0] operation_274_2658;
wire signed [31:0] operation_274_2657;
wire signed [31:0] operation_274_2656;
wire signed [31:0] operation_274_2655;
wire signed [31:0] operation_274_2654;
wire signed [31:0] operation_274_2653;
wire signed [31:0] operation_274_2652;
wire signed [31:0] operation_274_2651;
wire signed [31:0] operation_274_2650;
wire signed [31:0] operation_274_2649;
wire signed [31:0] operation_274_2648;
wire signed [31:0] operation_274_2647;
wire signed [31:0] operation_274_2646;
wire signed [31:0] operation_274_2645;
wire signed [31:0] operation_274_2644;
wire signed [31:0] operation_274_2643;
wire [7:0] operation_274_3109;
wire [7:0] operation_274_3108;
wire [7:0] operation_274_3090;
wire [7:0] operation_274_3036;
wire [7:0] operation_274_2678;
wire [7:0] operation_274_2677;
wire [7:0] operation_274_2676;
wire [7:0] operation_274_2675;
wire [7:0] operation_274_2674;
wire [7:0] operation_274_2673;
wire [7:0] operation_274_2672;
wire [7:0] operation_274_2671;
wire [7:0] operation_274_2670;
wire [7:0] operation_274_2669;
wire [7:0] operation_274_2668;
wire [7:0] operation_274_2667;
wire [7:0] operation_274_2666;
wire [7:0] operation_274_2665;
wire [7:0] operation_274_2664;
wire [7:0] operation_274_2663;
reg signed [31:0] operation_274_3129;
reg signed [31:0] operation_274_3128;
reg signed [31:0] operation_274_3110;
reg signed [31:0] operation_274_3053;
reg signed [31:0] operation_274_2698;
reg signed [31:0] operation_274_2697;
reg signed [31:0] operation_274_2696;
reg signed [31:0] operation_274_2695;
reg signed [31:0] operation_274_2694;
reg signed [31:0] operation_274_2693;
reg signed [31:0] operation_274_2692;
reg signed [31:0] operation_274_2691;
reg signed [31:0] operation_274_2690;
reg signed [31:0] operation_274_2689;
reg signed [31:0] operation_274_2688;
reg signed [31:0] operation_274_2687;
reg signed [31:0] operation_274_2686;
reg signed [31:0] operation_274_2685;
reg signed [31:0] operation_274_2684;
reg signed [31:0] operation_274_2683;
wire signed [31:0] operation_274_3149;
wire signed [31:0] operation_274_3148;
wire signed [31:0] operation_274_3130;
wire signed [31:0] operation_274_3071;
wire signed [31:0] operation_274_2718;
wire signed [31:0] operation_274_2717;
wire signed [31:0] operation_274_2716;
wire signed [31:0] operation_274_2715;
wire signed [31:0] operation_274_2714;
wire signed [31:0] operation_274_2713;
wire signed [31:0] operation_274_2712;
wire signed [31:0] operation_274_2711;
wire signed [31:0] operation_274_2710;
wire signed [31:0] operation_274_2709;
wire signed [31:0] operation_274_2708;
wire signed [31:0] operation_274_2707;
wire signed [31:0] operation_274_2706;
wire signed [31:0] operation_274_2705;
wire signed [31:0] operation_274_2704;
wire signed [31:0] operation_274_2703;
wire [7:0] operation_274_3169;
wire [7:0] operation_274_3168;
wire [7:0] operation_274_3150;
wire [7:0] operation_274_3091;
wire [7:0] operation_274_2738;
wire [7:0] operation_274_2737;
wire [7:0] operation_274_2736;
wire [7:0] operation_274_2735;
wire [7:0] operation_274_2734;
wire [7:0] operation_274_2733;
wire [7:0] operation_274_2732;
wire [7:0] operation_274_2731;
wire [7:0] operation_274_2730;
wire [7:0] operation_274_2729;
wire [7:0] operation_274_2728;
wire [7:0] operation_274_2727;
wire [7:0] operation_274_2726;
wire [7:0] operation_274_2725;
wire [7:0] operation_274_2724;
wire [7:0] operation_274_2723;
reg signed [31:0] operation_274_3189;
reg signed [31:0] operation_274_3188;
reg signed [31:0] operation_274_3170;
reg signed [31:0] operation_274_3111;
reg signed [31:0] operation_274_2758;
reg signed [31:0] operation_274_2757;
reg signed [31:0] operation_274_2756;
reg signed [31:0] operation_274_2755;
reg signed [31:0] operation_274_2754;
reg signed [31:0] operation_274_2753;
reg signed [31:0] operation_274_2752;
reg signed [31:0] operation_274_2751;
reg signed [31:0] operation_274_2750;
reg signed [31:0] operation_274_2749;
reg signed [31:0] operation_274_2748;
reg signed [31:0] operation_274_2747;
reg signed [31:0] operation_274_2746;
reg signed [31:0] operation_274_2745;
reg signed [31:0] operation_274_2744;
reg signed [31:0] operation_274_2743;
wire signed [31:0] operation_274_3209;
wire signed [31:0] operation_274_3208;
wire signed [31:0] operation_274_3190;
wire signed [31:0] operation_274_3131;
reg signed [31:0] operation_274_2778;
reg signed [31:0] operation_274_2777;
reg signed [31:0] operation_274_2776;
reg signed [31:0] operation_274_2775;
reg signed [31:0] operation_274_2774;
reg signed [31:0] operation_274_2773;
reg signed [31:0] operation_274_2772;
reg signed [31:0] operation_274_2771;
reg signed [31:0] operation_274_2770;
reg signed [31:0] operation_274_2769;
reg signed [31:0] operation_274_2768;
reg signed [31:0] operation_274_2767;
reg signed [31:0] operation_274_2766;
reg signed [31:0] operation_274_2765;
reg signed [31:0] operation_274_2764;
reg signed [31:0] operation_274_2763;
wire [7:0] operation_274_3233;
wire [7:0] operation_274_3232;
wire [7:0] operation_274_3210;
wire [7:0] operation_274_3151;
reg signed [31:0] operation_274_2802;
reg signed [31:0] operation_274_2801;
reg signed [31:0] operation_274_2800;
reg signed [31:0] operation_274_2799;
reg signed [31:0] operation_274_2798;
reg signed [31:0] operation_274_2797;
reg signed [31:0] operation_274_2796;
reg signed [31:0] operation_274_2795;
reg signed [31:0] operation_274_2794;
reg signed [31:0] operation_274_2793;
reg signed [31:0] operation_274_2792;
reg signed [31:0] operation_274_2791;
reg signed [31:0] operation_274_2790;
reg signed [31:0] operation_274_2789;
reg signed [31:0] operation_274_2788;
reg signed [31:0] operation_274_2787;
wire signed [31:0] operation_274_2786;
wire signed [31:0] operation_274_2785;
wire signed [31:0] operation_274_2784;
wire signed [31:0] operation_274_2783;
reg signed [31:0] operation_274_3273;
reg signed [31:0] operation_274_3272;
reg signed [31:0] operation_274_3234;
reg signed [31:0] operation_274_3171;
wire [7:0] operation_274_2842;
wire [7:0] operation_274_2841;
reg signed [31:0] operation_274_2840;
reg signed [31:0] operation_274_2839;
reg signed [31:0] operation_274_2838;
reg signed [31:0] operation_274_2837;
reg signed [31:0] operation_274_2836;
reg signed [31:0] operation_274_2835;
reg signed [31:0] operation_274_2834;
reg signed [31:0] operation_274_2833;
reg signed [31:0] operation_274_2832;
reg signed [31:0] operation_274_2831;
reg signed [31:0] operation_274_2830;
reg signed [31:0] operation_274_2829;
reg signed [31:0] operation_274_2828;
reg signed [31:0] operation_274_2827;
reg signed [31:0] operation_274_2826;
reg signed [31:0] operation_274_2825;
reg signed [31:0] operation_274_2824;
reg signed [31:0] operation_274_2823;
reg signed [31:0] operation_274_2822;
reg signed [31:0] operation_274_2821;
reg signed [31:0] operation_274_2820;
reg signed [31:0] operation_274_2819;
reg signed [31:0] operation_274_2818;
reg signed [31:0] operation_274_2817;
reg signed [31:0] operation_274_2816;
reg signed [31:0] operation_274_2815;
reg signed [31:0] operation_274_2814;
reg signed [31:0] operation_274_2813;
reg signed [31:0] operation_274_2812;
reg signed [31:0] operation_274_2811;
reg signed [31:0] operation_274_2810;
reg signed [31:0] operation_274_2809;
wire [7:0] operation_274_2808;
wire [7:0] operation_274_2807;
wire signed [31:0] operation_274_3297;
wire signed [31:0] operation_274_3296;
wire signed [31:0] operation_274_3274;
wire signed [31:0] operation_274_3191;
reg signed [31:0] operation_274_2866;
reg signed [31:0] operation_274_2865;
wire signed [31:0] operation_274_2864;
wire signed [31:0] operation_274_2863;
wire signed [31:0] operation_274_2862;
wire signed [31:0] operation_274_2861;
wire signed [31:0] operation_274_2860;
wire signed [31:0] operation_274_2859;
wire signed [31:0] operation_274_2858;
wire signed [31:0] operation_274_2857;
wire signed [31:0] operation_274_2856;
wire signed [31:0] operation_274_2855;
wire signed [31:0] operation_274_2854;
wire signed [31:0] operation_274_2853;
wire signed [31:0] operation_274_2852;
wire signed [31:0] operation_274_2851;
wire signed [31:0] operation_274_2850;
wire signed [31:0] operation_274_2849;
reg signed [31:0] operation_274_2848;
reg signed [31:0] operation_274_2847;
wire [7:0] operation_274_3322;
wire [7:0] operation_274_3321;
wire [7:0] operation_274_3299;
wire [7:0] operation_274_3211;
reg signed [31:0] operation_274_2890;
reg signed [31:0] operation_274_2889;
wire [7:0] operation_274_2888;
wire [7:0] operation_274_2887;
wire [7:0] operation_274_2886;
wire [7:0] operation_274_2885;
wire [7:0] operation_274_2884;
wire [7:0] operation_274_2883;
wire [7:0] operation_274_2882;
wire [7:0] operation_274_2881;
wire [7:0] operation_274_2880;
wire [7:0] operation_274_2879;
wire [7:0] operation_274_2878;
wire [7:0] operation_274_2877;
wire [7:0] operation_274_2876;
wire [7:0] operation_274_2875;
wire [7:0] operation_274_2874;
wire [7:0] operation_274_2873;
reg signed [31:0] operation_274_2872;
reg signed [31:0] operation_274_2871;
reg signed [31:0] operation_274_3343;
reg signed [31:0] operation_274_3342;
reg signed [31:0] operation_274_3324;
reg signed [31:0] operation_274_3235;
reg signed [31:0] operation_274_2911;
reg signed [31:0] operation_274_2910;
reg signed [31:0] operation_274_2909;
reg signed [31:0] operation_274_2908;
reg signed [31:0] operation_274_2907;
reg signed [31:0] operation_274_2906;
reg signed [31:0] operation_274_2905;
reg signed [31:0] operation_274_2904;
reg signed [31:0] operation_274_2903;
reg signed [31:0] operation_274_2902;
reg signed [31:0] operation_274_2901;
reg signed [31:0] operation_274_2900;
reg signed [31:0] operation_274_2899;
reg signed [31:0] operation_274_2898;
reg signed [31:0] operation_274_2897;
reg signed [31:0] operation_274_2896;
wire signed [31:0] operation_274_3365;
wire signed [31:0] operation_274_3364;
wire signed [31:0] operation_274_3346;
wire signed [31:0] operation_274_3275;
wire signed [31:0] operation_274_2933;
wire signed [31:0] operation_274_2932;
wire signed [31:0] operation_274_2931;
wire signed [31:0] operation_274_2930;
wire signed [31:0] operation_274_2929;
wire signed [31:0] operation_274_2928;
wire signed [31:0] operation_274_2927;
wire signed [31:0] operation_274_2926;
wire signed [31:0] operation_274_2925;
wire signed [31:0] operation_274_2924;
wire signed [31:0] operation_274_2923;
wire signed [31:0] operation_274_2922;
wire signed [31:0] operation_274_2921;
wire signed [31:0] operation_274_2920;
wire signed [31:0] operation_274_2919;
wire signed [31:0] operation_274_2918;
wire signed [31:0] operation_274_2660;
wire signed [31:0] operation_274_2641;
wire signed [31:0] operation_274_2590;
reg [7:0] operation_274_3393_latch;
wire [7:0] operation_274_3393;
reg [7:0] operation_274_3375_latch;
wire [7:0] operation_274_3375;
reg [7:0] operation_274_3374_latch;
wire [7:0] operation_274_3374;
wire [7:0] operation_274_3320;
reg [7:0] operation_274_2962_latch;
wire [7:0] operation_274_2962;
reg [7:0] operation_274_2961_latch;
wire [7:0] operation_274_2961;
reg [7:0] operation_274_2960_latch;
wire [7:0] operation_274_2960;
reg [7:0] operation_274_2959_latch;
wire [7:0] operation_274_2959;
reg [7:0] operation_274_2958_latch;
wire [7:0] operation_274_2958;
reg [7:0] operation_274_2957_latch;
wire [7:0] operation_274_2957;
reg [7:0] operation_274_2956_latch;
wire [7:0] operation_274_2956;
reg [7:0] operation_274_2955_latch;
wire [7:0] operation_274_2955;
reg [7:0] operation_274_2954_latch;
wire [7:0] operation_274_2954;
reg [7:0] operation_274_2953_latch;
wire [7:0] operation_274_2953;
reg [7:0] operation_274_2952_latch;
wire [7:0] operation_274_2952;
reg [7:0] operation_274_2951_latch;
wire [7:0] operation_274_2951;
reg [7:0] operation_274_2950_latch;
wire [7:0] operation_274_2950;
reg [7:0] operation_274_2949_latch;
wire [7:0] operation_274_2949;
reg [7:0] operation_274_2948_latch;
wire [7:0] operation_274_2948;
reg [7:0] operation_274_2947_latch;
wire [7:0] operation_274_2947;
wire [7:0] operation_274_2680;
wire [7:0] operation_274_2661;
wire [7:0] operation_274_2607;
reg signed [31:0] operation_274_3341;
wire [7:0] operation_274_2143;
wire [7:0] operation_274_2142;
wire [7:0] operation_274_2141;
wire [7:0] operation_274_2140;
wire [7:0] operation_274_2139;
wire [7:0] operation_274_2138;
wire [7:0] operation_274_2137;
wire [7:0] operation_274_2136;
wire [7:0] operation_274_2135;
wire [7:0] operation_274_2134;
wire [7:0] operation_274_2133;
wire [7:0] operation_274_2132;
wire [7:0] operation_274_2131;
wire [7:0] operation_274_2130;
wire [7:0] operation_274_2129;
wire [7:0] operation_274_2128;
reg signed [31:0] operation_274_2700;
reg signed [31:0] operation_274_2681;
reg signed [31:0] operation_274_2624;
wire signed [31:0] operation_274_3363;
reg signed [31:0] operation_274_2159;
reg signed [31:0] operation_274_2158;
reg signed [31:0] operation_274_2157;
reg signed [31:0] operation_274_2156;
reg signed [31:0] operation_274_2155;
reg signed [31:0] operation_274_2154;
reg signed [31:0] operation_274_2153;
reg signed [31:0] operation_274_2152;
reg signed [31:0] operation_274_2151;
reg signed [31:0] operation_274_2150;
reg signed [31:0] operation_274_2149;
reg signed [31:0] operation_274_2148;
reg signed [31:0] operation_274_2147;
reg signed [31:0] operation_274_2146;
reg signed [31:0] operation_274_2145;
reg signed [31:0] operation_274_2144;
wire signed [31:0] operation_274_2720;
wire signed [31:0] operation_274_2701;
wire signed [31:0] operation_274_2659;
wire signed [31:0] operation_274_2642;
reg [7:0] operation_274_3392_latch;
wire [7:0] operation_274_3392;
wire signed [31:0] operation_274_2177;
wire signed [31:0] operation_274_2176;
wire signed [31:0] operation_274_2175;
wire signed [31:0] operation_274_2174;
wire signed [31:0] operation_274_2173;
wire signed [31:0] operation_274_2172;
wire signed [31:0] operation_274_2171;
wire signed [31:0] operation_274_2170;
wire signed [31:0] operation_274_2168;
wire signed [31:0] operation_274_2167;
wire signed [31:0] operation_274_2166;
wire signed [31:0] operation_274_2165;
wire signed [31:0] operation_274_2164;
wire signed [31:0] operation_274_2163;
wire signed [31:0] operation_274_2162;
wire signed [31:0] operation_274_2160;
wire [7:0] operation_274_2740;
wire [7:0] operation_274_2721;
wire [7:0] operation_274_2679;
wire [7:0] operation_274_2662;
wire [7:0] operation_274_2194;
wire [7:0] operation_274_2193;
wire [7:0] operation_274_2192;
wire [7:0] operation_274_2191;
wire [7:0] operation_274_2190;
wire [7:0] operation_274_2189;
wire [7:0] operation_274_2188;
wire [7:0] operation_274_2187;
wire [7:0] operation_274_2186;
wire [7:0] operation_274_2185;
wire [7:0] operation_274_2184;
wire [7:0] operation_274_2183;
wire [7:0] operation_274_2182;
wire [7:0] operation_274_2181;
wire [7:0] operation_274_2180;
wire [7:0] operation_274_2179;
reg signed [31:0] operation_274_2760;
reg signed [31:0] operation_274_2741;
reg signed [31:0] operation_274_2699;
reg signed [31:0] operation_274_2682;
reg signed [31:0] operation_274_2211;
reg signed [31:0] operation_274_2210;
reg signed [31:0] operation_274_2209;
reg signed [31:0] operation_274_2208;
reg signed [31:0] operation_274_2207;
reg signed [31:0] operation_274_2206;
reg signed [31:0] operation_274_2205;
reg signed [31:0] operation_274_2204;
reg signed [31:0] operation_274_2203;
reg signed [31:0] operation_274_2202;
reg signed [31:0] operation_274_2201;
reg signed [31:0] operation_274_2200;
reg signed [31:0] operation_274_2199;
reg signed [31:0] operation_274_2198;
reg signed [31:0] operation_274_2197;
reg signed [31:0] operation_274_2196;
wire signed [31:0] operation_274_2780;
wire signed [31:0] operation_274_2761;
wire signed [31:0] operation_274_2719;
wire signed [31:0] operation_274_2702;
wire signed [31:0] operation_274_2229;
wire signed [31:0] operation_274_2228;
wire signed [31:0] operation_274_2227;
wire signed [31:0] operation_274_2226;
wire signed [31:0] operation_274_2225;
wire signed [31:0] operation_274_2224;
wire signed [31:0] operation_274_2223;
wire signed [31:0] operation_274_2222;
wire signed [31:0] operation_274_2221;
wire signed [31:0] operation_274_2220;
wire signed [31:0] operation_274_2219;
wire signed [31:0] operation_274_2218;
wire signed [31:0] operation_274_2217;
wire signed [31:0] operation_274_2216;
wire signed [31:0] operation_274_2215;
wire signed [31:0] operation_274_2214;
wire [7:0] operation_274_2804;
wire [7:0] operation_274_2781;
wire [7:0] operation_274_2739;
wire [7:0] operation_274_2722;
wire [7:0] operation_274_2249;
wire [7:0] operation_274_2248;
wire [7:0] operation_274_2247;
wire [7:0] operation_274_2246;
wire [7:0] operation_274_2245;
wire [7:0] operation_274_2244;
wire [7:0] operation_274_2243;
wire [7:0] operation_274_2242;
wire [7:0] operation_274_2241;
wire [7:0] operation_274_2240;
wire [7:0] operation_274_2239;
wire [7:0] operation_274_2238;
wire [7:0] operation_274_2237;
wire [7:0] operation_274_2236;
wire [7:0] operation_274_2235;
wire [7:0] operation_274_2234;
reg signed [31:0] operation_274_2844;
reg signed [31:0] operation_274_2805;
reg signed [31:0] operation_274_2759;
reg signed [31:0] operation_274_2742;
reg signed [31:0] operation_274_2269;
reg signed [31:0] operation_274_2268;
reg signed [31:0] operation_274_2267;
reg signed [31:0] operation_274_2266;
reg signed [31:0] operation_274_2265;
reg signed [31:0] operation_274_2264;
reg signed [31:0] operation_274_2263;
reg signed [31:0] operation_274_2262;
reg signed [31:0] operation_274_2261;
reg signed [31:0] operation_274_2260;
reg signed [31:0] operation_274_2259;
reg signed [31:0] operation_274_2258;
reg signed [31:0] operation_274_2257;
reg signed [31:0] operation_274_2256;
reg signed [31:0] operation_274_2255;
reg signed [31:0] operation_274_2254;
wire signed [31:0] operation_274_2868;
wire signed [31:0] operation_274_2845;
wire signed [31:0] operation_274_2779;
wire signed [31:0] operation_274_2762;
wire signed [31:0] operation_274_2289;
wire signed [31:0] operation_274_2288;
wire signed [31:0] operation_274_2287;
wire signed [31:0] operation_274_2286;
wire signed [31:0] operation_274_2285;
wire signed [31:0] operation_274_2284;
wire signed [31:0] operation_274_2283;
wire signed [31:0] operation_274_2282;
wire signed [31:0] operation_274_2281;
wire signed [31:0] operation_274_2280;
wire signed [31:0] operation_274_2279;
wire signed [31:0] operation_274_2278;
wire signed [31:0] operation_274_2277;
wire signed [31:0] operation_274_2276;
wire signed [31:0] operation_274_2275;
wire signed [31:0] operation_274_2274;
wire [7:0] operation_274_2893;
wire [7:0] operation_274_2870;
wire [7:0] operation_274_2803;
wire [7:0] operation_274_2782;
wire [7:0] operation_274_2309;
wire [7:0] operation_274_2308;
wire [7:0] operation_274_2307;
wire [7:0] operation_274_2306;
wire [7:0] operation_274_2305;
wire [7:0] operation_274_2304;
wire [7:0] operation_274_2303;
wire [7:0] operation_274_2302;
wire [7:0] operation_274_2301;
wire [7:0] operation_274_2300;
wire [7:0] operation_274_2299;
wire [7:0] operation_274_2298;
wire [7:0] operation_274_2297;
wire [7:0] operation_274_2296;
wire [7:0] operation_274_2295;
wire [7:0] operation_274_2294;
reg signed [31:0] operation_274_2914;
reg signed [31:0] operation_274_2895;
reg signed [31:0] operation_274_2843;
reg signed [31:0] operation_274_2806;
reg signed [31:0] operation_274_2329;
reg signed [31:0] operation_274_2328;
reg signed [31:0] operation_274_2327;
reg signed [31:0] operation_274_2326;
reg signed [31:0] operation_274_2325;
reg signed [31:0] operation_274_2324;
reg signed [31:0] operation_274_2323;
reg signed [31:0] operation_274_2322;
reg signed [31:0] operation_274_2321;
reg signed [31:0] operation_274_2320;
reg signed [31:0] operation_274_2319;
reg signed [31:0] operation_274_2318;
reg signed [31:0] operation_274_2317;
reg signed [31:0] operation_274_2316;
reg signed [31:0] operation_274_2315;
reg signed [31:0] operation_274_2314;
wire signed [31:0] operation_274_2936;
wire signed [31:0] operation_274_2917;
wire signed [31:0] operation_274_2867;
wire signed [31:0] operation_274_2846;
reg signed [31:0] operation_274_2349;
reg signed [31:0] operation_274_2348;
reg signed [31:0] operation_274_2347;
reg signed [31:0] operation_274_2346;
reg signed [31:0] operation_274_2345;
reg signed [31:0] operation_274_2344;
reg signed [31:0] operation_274_2343;
reg signed [31:0] operation_274_2342;
reg signed [31:0] operation_274_2341;
reg signed [31:0] operation_274_2340;
reg signed [31:0] operation_274_2339;
reg signed [31:0] operation_274_2338;
reg signed [31:0] operation_274_2337;
reg signed [31:0] operation_274_2336;
reg signed [31:0] operation_274_2335;
reg signed [31:0] operation_274_2334;
wire signed [31:0] operation_274_2231;
wire signed [31:0] operation_274_2161;
reg [7:0] operation_274_2964_latch;
wire [7:0] operation_274_2964;
reg [7:0] operation_274_2945_latch;
wire [7:0] operation_274_2945;
wire [7:0] operation_274_2892;
wire [7:0] operation_274_2891;
reg signed [31:0] operation_274_2373;
reg signed [31:0] operation_274_2372;
reg signed [31:0] operation_274_2371;
reg signed [31:0] operation_274_2370;
reg signed [31:0] operation_274_2369;
reg signed [31:0] operation_274_2368;
reg signed [31:0] operation_274_2367;
reg signed [31:0] operation_274_2366;
reg signed [31:0] operation_274_2365;
reg signed [31:0] operation_274_2364;
reg signed [31:0] operation_274_2363;
reg signed [31:0] operation_274_2362;
reg signed [31:0] operation_274_2361;
reg signed [31:0] operation_274_2360;
reg signed [31:0] operation_274_2359;
reg signed [31:0] operation_274_2358;
wire signed [31:0] operation_274_2357;
wire signed [31:0] operation_274_2356;
wire signed [31:0] operation_274_2355;
wire signed [31:0] operation_274_2354;
wire [7:0] operation_274_2251;
wire [7:0] operation_274_2178;
reg signed [31:0] operation_274_2913;
reg signed [31:0] operation_274_2912;
wire [7:0] operation_274_2413;
wire [7:0] operation_274_2412;
reg signed [31:0] operation_274_2411;
reg signed [31:0] operation_274_2410;
reg signed [31:0] operation_274_2409;
reg signed [31:0] operation_274_2408;
reg signed [31:0] operation_274_2407;
reg signed [31:0] operation_274_2406;
reg signed [31:0] operation_274_2405;
reg signed [31:0] operation_274_2404;
reg signed [31:0] operation_274_2403;
reg signed [31:0] operation_274_2402;
reg signed [31:0] operation_274_2401;
reg signed [31:0] operation_274_2400;
reg signed [31:0] operation_274_2399;
reg signed [31:0] operation_274_2398;
reg signed [31:0] operation_274_2397;
reg signed [31:0] operation_274_2396;
reg signed [31:0] operation_274_2395;
reg signed [31:0] operation_274_2394;
reg signed [31:0] operation_274_2393;
reg signed [31:0] operation_274_2392;
reg signed [31:0] operation_274_2391;
reg signed [31:0] operation_274_2390;
reg signed [31:0] operation_274_2389;
reg signed [31:0] operation_274_2388;
reg signed [31:0] operation_274_2387;
reg signed [31:0] operation_274_2386;
reg signed [31:0] operation_274_2385;
reg signed [31:0] operation_274_2384;
reg signed [31:0] operation_274_2383;
reg signed [31:0] operation_274_2382;
reg signed [31:0] operation_274_2381;
reg signed [31:0] operation_274_2380;
wire [7:0] operation_274_2379;
wire [7:0] operation_274_2378;
reg signed [31:0] operation_274_2271;
reg signed [31:0] operation_274_2195;
wire signed [31:0] operation_274_2935;
wire signed [31:0] operation_274_2934;
reg signed [31:0] operation_274_2437;
reg signed [31:0] operation_274_2436;
wire signed [31:0] operation_274_2435;
wire signed [31:0] operation_274_2434;
wire signed [31:0] operation_274_2433;
wire signed [31:0] operation_274_2432;
wire signed [31:0] operation_274_2431;
wire signed [31:0] operation_274_2430;
wire signed [31:0] operation_274_2429;
wire signed [31:0] operation_274_2428;
wire signed [31:0] operation_274_2427;
wire signed [31:0] operation_274_2426;
wire signed [31:0] operation_274_2425;
wire signed [31:0] operation_274_2424;
wire signed [31:0] operation_274_2423;
wire signed [31:0] operation_274_2422;
wire signed [31:0] operation_274_2421;
wire signed [31:0] operation_274_2420;
reg signed [31:0] operation_274_2419;
reg signed [31:0] operation_274_2418;
wire signed [31:0] operation_274_2291;
wire signed [31:0] operation_274_2230;
wire signed [31:0] operation_274_2213;
wire signed [31:0] operation_274_2212;
reg [7:0] operation_274_2963_latch;
wire [7:0] operation_274_2963;
reg [7:0] operation_274_2946_latch;
wire [7:0] operation_274_2946;
reg signed [31:0] operation_274_2461;
reg signed [31:0] operation_274_2460;
wire [7:0] operation_274_2459;
wire [7:0] operation_274_2458;
wire [7:0] operation_274_2457;
wire [7:0] operation_274_2456;
wire [7:0] operation_274_2455;
wire [7:0] operation_274_2454;
wire [7:0] operation_274_2453;
wire [7:0] operation_274_2452;
wire [7:0] operation_274_2451;
wire [7:0] operation_274_2450;
wire [7:0] operation_274_2449;
wire [7:0] operation_274_2448;
wire [7:0] operation_274_2447;
wire [7:0] operation_274_2446;
wire [7:0] operation_274_2445;
wire [7:0] operation_274_2444;
reg signed [31:0] operation_274_2443;
reg signed [31:0] operation_274_2442;
wire [7:0] operation_274_2311;
wire [7:0] operation_274_2250;
wire [7:0] operation_274_2233;
wire [7:0] operation_274_2232;
reg signed [31:0] operation_274_2482;
reg signed [31:0] operation_274_2481;
reg signed [31:0] operation_274_2480;
reg signed [31:0] operation_274_2479;
reg signed [31:0] operation_274_2478;
reg signed [31:0] operation_274_2477;
reg signed [31:0] operation_274_2476;
reg signed [31:0] operation_274_2475;
reg signed [31:0] operation_274_2474;
reg signed [31:0] operation_274_2473;
reg signed [31:0] operation_274_2472;
reg signed [31:0] operation_274_2471;
reg signed [31:0] operation_274_2470;
reg signed [31:0] operation_274_2469;
reg signed [31:0] operation_274_2468;
reg signed [31:0] operation_274_2467;
reg signed [31:0] operation_274_2331;
reg signed [31:0] operation_274_2270;
reg signed [31:0] operation_274_2253;
reg signed [31:0] operation_274_2252;
wire signed [31:0] operation_274_2504;
wire signed [31:0] operation_274_2503;
wire signed [31:0] operation_274_2502;
wire signed [31:0] operation_274_2501;
wire signed [31:0] operation_274_2500;
wire signed [31:0] operation_274_2499;
wire signed [31:0] operation_274_2498;
wire signed [31:0] operation_274_2497;
wire signed [31:0] operation_274_2496;
wire signed [31:0] operation_274_2495;
wire signed [31:0] operation_274_2494;
wire signed [31:0] operation_274_2493;
wire signed [31:0] operation_274_2492;
wire signed [31:0] operation_274_2491;
wire signed [31:0] operation_274_2490;
wire signed [31:0] operation_274_2489;
wire signed [31:0] operation_274_2351;
wire signed [31:0] operation_274_2290;
wire signed [31:0] operation_274_2273;
wire signed [31:0] operation_274_2272;
reg [7:0] operation_274_2533_latch;
wire [7:0] operation_274_2533;
reg [7:0] operation_274_2532_latch;
wire [7:0] operation_274_2532;
reg [7:0] operation_274_2531_latch;
wire [7:0] operation_274_2531;
reg [7:0] operation_274_2530_latch;
wire [7:0] operation_274_2530;
reg [7:0] operation_274_2529_latch;
wire [7:0] operation_274_2529;
reg [7:0] operation_274_2528_latch;
wire [7:0] operation_274_2528;
reg [7:0] operation_274_2527_latch;
wire [7:0] operation_274_2527;
reg [7:0] operation_274_2526_latch;
wire [7:0] operation_274_2526;
reg [7:0] operation_274_2525_latch;
wire [7:0] operation_274_2525;
reg [7:0] operation_274_2524_latch;
wire [7:0] operation_274_2524;
reg [7:0] operation_274_2523_latch;
wire [7:0] operation_274_2523;
reg [7:0] operation_274_2522_latch;
wire [7:0] operation_274_2522;
reg [7:0] operation_274_2521_latch;
wire [7:0] operation_274_2521;
reg [7:0] operation_274_2520_latch;
wire [7:0] operation_274_2520;
reg [7:0] operation_274_2519_latch;
wire [7:0] operation_274_2519;
reg [7:0] operation_274_2518_latch;
wire [7:0] operation_274_2518;
wire [7:0] operation_274_2375;
wire [7:0] operation_274_2310;
wire [7:0] operation_274_2293;
wire [7:0] operation_274_2292;
wire [7:0] operation_274_1714;
wire [7:0] operation_274_1713;
wire [7:0] operation_274_1712;
wire [7:0] operation_274_1711;
wire [7:0] operation_274_1710;
wire [7:0] operation_274_1709;
wire [7:0] operation_274_1708;
wire [7:0] operation_274_1707;
wire [7:0] operation_274_1706;
wire [7:0] operation_274_1705;
wire [7:0] operation_274_1704;
wire [7:0] operation_274_1703;
wire [7:0] operation_274_1702;
wire [7:0] operation_274_1701;
wire [7:0] operation_274_1700;
wire [7:0] operation_274_1699;
reg signed [31:0] operation_274_2415;
reg signed [31:0] operation_274_2330;
reg signed [31:0] operation_274_2313;
reg signed [31:0] operation_274_2312;
reg signed [31:0] operation_274_1730;
reg signed [31:0] operation_274_1729;
reg signed [31:0] operation_274_1728;
reg signed [31:0] operation_274_1727;
reg signed [31:0] operation_274_1726;
reg signed [31:0] operation_274_1725;
reg signed [31:0] operation_274_1724;
reg signed [31:0] operation_274_1723;
reg signed [31:0] operation_274_1722;
reg signed [31:0] operation_274_1721;
reg signed [31:0] operation_274_1720;
reg signed [31:0] operation_274_1719;
reg signed [31:0] operation_274_1718;
reg signed [31:0] operation_274_1717;
reg signed [31:0] operation_274_1716;
reg signed [31:0] operation_274_1715;
wire signed [31:0] operation_274_2439;
wire signed [31:0] operation_274_2350;
wire signed [31:0] operation_274_2333;
wire signed [31:0] operation_274_2332;
wire signed [31:0] operation_274_1748;
wire signed [31:0] operation_274_1747;
wire signed [31:0] operation_274_1746;
wire signed [31:0] operation_274_1745;
wire signed [31:0] operation_274_1744;
wire signed [31:0] operation_274_1743;
wire signed [31:0] operation_274_1742;
wire signed [31:0] operation_274_1741;
wire signed [31:0] operation_274_1739;
wire signed [31:0] operation_274_1738;
wire signed [31:0] operation_274_1737;
wire signed [31:0] operation_274_1736;
wire signed [31:0] operation_274_1735;
wire signed [31:0] operation_274_1734;
wire signed [31:0] operation_274_1733;
wire signed [31:0] operation_274_1731;
wire [7:0] operation_274_2464;
wire [7:0] operation_274_2374;
wire [7:0] operation_274_2353;
wire [7:0] operation_274_2352;
wire [7:0] operation_274_1765;
wire [7:0] operation_274_1764;
wire [7:0] operation_274_1763;
wire [7:0] operation_274_1762;
wire [7:0] operation_274_1761;
wire [7:0] operation_274_1760;
wire [7:0] operation_274_1759;
wire [7:0] operation_274_1758;
wire [7:0] operation_274_1757;
wire [7:0] operation_274_1756;
wire [7:0] operation_274_1755;
wire [7:0] operation_274_1754;
wire [7:0] operation_274_1753;
wire [7:0] operation_274_1752;
wire [7:0] operation_274_1751;
wire [7:0] operation_274_1750;
reg signed [31:0] operation_274_2485;
reg signed [31:0] operation_274_2414;
reg signed [31:0] operation_274_2377;
reg signed [31:0] operation_274_2376;
reg signed [31:0] operation_274_1782;
reg signed [31:0] operation_274_1781;
reg signed [31:0] operation_274_1780;
reg signed [31:0] operation_274_1779;
reg signed [31:0] operation_274_1778;
reg signed [31:0] operation_274_1777;
reg signed [31:0] operation_274_1776;
reg signed [31:0] operation_274_1775;
reg signed [31:0] operation_274_1774;
reg signed [31:0] operation_274_1773;
reg signed [31:0] operation_274_1772;
reg signed [31:0] operation_274_1771;
reg signed [31:0] operation_274_1770;
reg signed [31:0] operation_274_1769;
reg signed [31:0] operation_274_1768;
reg signed [31:0] operation_274_1767;
wire signed [31:0] operation_274_2507;
wire signed [31:0] operation_274_2438;
wire signed [31:0] operation_274_2417;
wire signed [31:0] operation_274_2416;
wire signed [31:0] operation_274_1800;
wire signed [31:0] operation_274_1799;
wire signed [31:0] operation_274_1798;
wire signed [31:0] operation_274_1797;
wire signed [31:0] operation_274_1796;
wire signed [31:0] operation_274_1795;
wire signed [31:0] operation_274_1794;
wire signed [31:0] operation_274_1793;
wire signed [31:0] operation_274_1792;
wire signed [31:0] operation_274_1791;
wire signed [31:0] operation_274_1790;
wire signed [31:0] operation_274_1789;
wire signed [31:0] operation_274_1788;
wire signed [31:0] operation_274_1787;
wire signed [31:0] operation_274_1786;
wire signed [31:0] operation_274_1785;
wire signed [31:0] operation_274_1732;
reg [7:0] operation_274_2516_latch;
wire [7:0] operation_274_2516;
wire [7:0] operation_274_2463;
wire [7:0] operation_274_2462;
wire [7:0] operation_274_2441;
wire [7:0] operation_274_1820;
wire [7:0] operation_274_1819;
wire [7:0] operation_274_1818;
wire [7:0] operation_274_1817;
wire [7:0] operation_274_1816;
wire [7:0] operation_274_1815;
wire [7:0] operation_274_1814;
wire [7:0] operation_274_1813;
wire [7:0] operation_274_1812;
wire [7:0] operation_274_1811;
wire [7:0] operation_274_1810;
wire [7:0] operation_274_1809;
wire [7:0] operation_274_1808;
wire [7:0] operation_274_1807;
wire [7:0] operation_274_1806;
wire [7:0] operation_274_1805;
wire [7:0] operation_274_1749;
reg signed [31:0] operation_274_2484;
reg signed [31:0] operation_274_2483;
reg signed [31:0] operation_274_2466;
reg signed [31:0] operation_274_1840;
reg signed [31:0] operation_274_1839;
reg signed [31:0] operation_274_1838;
reg signed [31:0] operation_274_1837;
reg signed [31:0] operation_274_1836;
reg signed [31:0] operation_274_1835;
reg signed [31:0] operation_274_1834;
reg signed [31:0] operation_274_1833;
reg signed [31:0] operation_274_1832;
reg signed [31:0] operation_274_1831;
reg signed [31:0] operation_274_1830;
reg signed [31:0] operation_274_1829;
reg signed [31:0] operation_274_1828;
reg signed [31:0] operation_274_1827;
reg signed [31:0] operation_274_1826;
reg signed [31:0] operation_274_1825;
reg signed [31:0] operation_274_1766;
wire signed [31:0] operation_274_2506;
wire signed [31:0] operation_274_2505;
wire signed [31:0] operation_274_2488;
wire signed [31:0] operation_274_1860;
wire signed [31:0] operation_274_1859;
wire signed [31:0] operation_274_1858;
wire signed [31:0] operation_274_1857;
wire signed [31:0] operation_274_1856;
wire signed [31:0] operation_274_1855;
wire signed [31:0] operation_274_1854;
wire signed [31:0] operation_274_1853;
wire signed [31:0] operation_274_1852;
wire signed [31:0] operation_274_1851;
wire signed [31:0] operation_274_1850;
wire signed [31:0] operation_274_1849;
wire signed [31:0] operation_274_1848;
wire signed [31:0] operation_274_1847;
wire signed [31:0] operation_274_1846;
wire signed [31:0] operation_274_1845;
wire signed [31:0] operation_274_1802;
wire signed [31:0] operation_274_1801;
wire signed [31:0] operation_274_1784;
wire signed [31:0] operation_274_1783;
reg [7:0] operation_274_2535_latch;
wire [7:0] operation_274_2535;
reg [7:0] operation_274_2534_latch;
wire [7:0] operation_274_2534;
reg [7:0] operation_274_2517_latch;
wire [7:0] operation_274_2517;
wire [7:0] operation_274_1880;
wire [7:0] operation_274_1879;
wire [7:0] operation_274_1878;
wire [7:0] operation_274_1877;
wire [7:0] operation_274_1876;
wire [7:0] operation_274_1875;
wire [7:0] operation_274_1874;
wire [7:0] operation_274_1873;
wire [7:0] operation_274_1872;
wire [7:0] operation_274_1871;
wire [7:0] operation_274_1870;
wire [7:0] operation_274_1869;
wire [7:0] operation_274_1868;
wire [7:0] operation_274_1867;
wire [7:0] operation_274_1866;
wire [7:0] operation_274_1865;
wire [7:0] operation_274_1822;
wire [7:0] operation_274_1821;
wire [7:0] operation_274_1804;
wire [7:0] operation_274_1803;
reg signed [31:0] operation_274_1900;
reg signed [31:0] operation_274_1899;
reg signed [31:0] operation_274_1898;
reg signed [31:0] operation_274_1897;
reg signed [31:0] operation_274_1896;
reg signed [31:0] operation_274_1895;
reg signed [31:0] operation_274_1894;
reg signed [31:0] operation_274_1893;
reg signed [31:0] operation_274_1892;
reg signed [31:0] operation_274_1891;
reg signed [31:0] operation_274_1890;
reg signed [31:0] operation_274_1889;
reg signed [31:0] operation_274_1888;
reg signed [31:0] operation_274_1887;
reg signed [31:0] operation_274_1886;
reg signed [31:0] operation_274_1885;
reg signed [31:0] operation_274_1842;
reg signed [31:0] operation_274_1841;
reg signed [31:0] operation_274_1824;
reg signed [31:0] operation_274_1823;
reg signed [31:0] operation_274_1920;
reg signed [31:0] operation_274_1919;
reg signed [31:0] operation_274_1918;
reg signed [31:0] operation_274_1917;
reg signed [31:0] operation_274_1916;
reg signed [31:0] operation_274_1915;
reg signed [31:0] operation_274_1914;
reg signed [31:0] operation_274_1913;
reg signed [31:0] operation_274_1912;
reg signed [31:0] operation_274_1911;
reg signed [31:0] operation_274_1910;
reg signed [31:0] operation_274_1909;
reg signed [31:0] operation_274_1908;
reg signed [31:0] operation_274_1907;
reg signed [31:0] operation_274_1906;
reg signed [31:0] operation_274_1905;
wire signed [31:0] operation_274_1862;
wire signed [31:0] operation_274_1861;
wire signed [31:0] operation_274_1844;
wire signed [31:0] operation_274_1843;
reg signed [31:0] operation_274_1944;
reg signed [31:0] operation_274_1943;
reg signed [31:0] operation_274_1942;
reg signed [31:0] operation_274_1941;
reg signed [31:0] operation_274_1940;
reg signed [31:0] operation_274_1939;
reg signed [31:0] operation_274_1938;
reg signed [31:0] operation_274_1937;
reg signed [31:0] operation_274_1936;
reg signed [31:0] operation_274_1935;
reg signed [31:0] operation_274_1934;
reg signed [31:0] operation_274_1933;
reg signed [31:0] operation_274_1932;
reg signed [31:0] operation_274_1931;
reg signed [31:0] operation_274_1930;
reg signed [31:0] operation_274_1929;
wire signed [31:0] operation_274_1928;
wire signed [31:0] operation_274_1927;
wire signed [31:0] operation_274_1926;
wire signed [31:0] operation_274_1925;
wire [7:0] operation_274_1882;
wire [7:0] operation_274_1881;
wire [7:0] operation_274_1864;
wire [7:0] operation_274_1863;
wire [7:0] operation_274_1984;
wire [7:0] operation_274_1983;
reg signed [31:0] operation_274_1982;
reg signed [31:0] operation_274_1981;
reg signed [31:0] operation_274_1980;
reg signed [31:0] operation_274_1979;
reg signed [31:0] operation_274_1978;
reg signed [31:0] operation_274_1977;
reg signed [31:0] operation_274_1976;
reg signed [31:0] operation_274_1975;
reg signed [31:0] operation_274_1974;
reg signed [31:0] operation_274_1973;
reg signed [31:0] operation_274_1972;
reg signed [31:0] operation_274_1971;
reg signed [31:0] operation_274_1970;
reg signed [31:0] operation_274_1969;
reg signed [31:0] operation_274_1968;
reg signed [31:0] operation_274_1967;
reg signed [31:0] operation_274_1966;
reg signed [31:0] operation_274_1965;
reg signed [31:0] operation_274_1964;
reg signed [31:0] operation_274_1963;
reg signed [31:0] operation_274_1962;
reg signed [31:0] operation_274_1961;
reg signed [31:0] operation_274_1960;
reg signed [31:0] operation_274_1959;
reg signed [31:0] operation_274_1958;
reg signed [31:0] operation_274_1957;
reg signed [31:0] operation_274_1956;
reg signed [31:0] operation_274_1955;
reg signed [31:0] operation_274_1954;
reg signed [31:0] operation_274_1953;
reg signed [31:0] operation_274_1952;
reg signed [31:0] operation_274_1951;
wire [7:0] operation_274_1950;
wire [7:0] operation_274_1949;
reg signed [31:0] operation_274_1902;
reg signed [31:0] operation_274_1901;
reg signed [31:0] operation_274_1884;
reg signed [31:0] operation_274_1883;
reg signed [31:0] operation_274_2008;
reg signed [31:0] operation_274_2007;
wire signed [31:0] operation_274_2006;
wire signed [31:0] operation_274_2005;
wire signed [31:0] operation_274_2004;
wire signed [31:0] operation_274_2003;
wire signed [31:0] operation_274_2002;
wire signed [31:0] operation_274_2001;
wire signed [31:0] operation_274_2000;
wire signed [31:0] operation_274_1999;
wire signed [31:0] operation_274_1998;
wire signed [31:0] operation_274_1997;
wire signed [31:0] operation_274_1996;
wire signed [31:0] operation_274_1995;
wire signed [31:0] operation_274_1994;
wire signed [31:0] operation_274_1993;
wire signed [31:0] operation_274_1992;
wire signed [31:0] operation_274_1991;
reg signed [31:0] operation_274_1990;
reg signed [31:0] operation_274_1989;
wire signed [31:0] operation_274_1922;
wire signed [31:0] operation_274_1921;
wire signed [31:0] operation_274_1904;
wire signed [31:0] operation_274_1903;
reg signed [31:0] operation_274_2032;
reg signed [31:0] operation_274_2031;
wire [7:0] operation_274_2030;
wire [7:0] operation_274_2029;
wire [7:0] operation_274_2028;
wire [7:0] operation_274_2027;
wire [7:0] operation_274_2026;
wire [7:0] operation_274_2025;
wire [7:0] operation_274_2024;
wire [7:0] operation_274_2023;
wire [7:0] operation_274_2022;
wire [7:0] operation_274_2021;
wire [7:0] operation_274_2020;
wire [7:0] operation_274_2019;
wire [7:0] operation_274_2018;
wire [7:0] operation_274_2017;
wire [7:0] operation_274_2016;
wire [7:0] operation_274_2015;
reg signed [31:0] operation_274_2014;
reg signed [31:0] operation_274_2013;
wire [7:0] operation_274_1946;
wire [7:0] operation_274_1945;
wire [7:0] operation_274_1924;
wire [7:0] operation_274_1923;
reg signed [31:0] operation_274_2053;
reg signed [31:0] operation_274_2052;
reg signed [31:0] operation_274_2051;
reg signed [31:0] operation_274_2050;
reg signed [31:0] operation_274_2049;
reg signed [31:0] operation_274_2048;
reg signed [31:0] operation_274_2047;
reg signed [31:0] operation_274_2046;
reg signed [31:0] operation_274_2045;
reg signed [31:0] operation_274_2044;
reg signed [31:0] operation_274_2043;
reg signed [31:0] operation_274_2042;
reg signed [31:0] operation_274_2041;
reg signed [31:0] operation_274_2040;
reg signed [31:0] operation_274_2039;
reg signed [31:0] operation_274_2038;
reg signed [31:0] operation_274_1986;
reg signed [31:0] operation_274_1985;
reg signed [31:0] operation_274_1948;
reg signed [31:0] operation_274_1947;
wire signed [31:0] operation_274_2075;
wire signed [31:0] operation_274_2074;
wire signed [31:0] operation_274_2073;
wire signed [31:0] operation_274_2072;
wire signed [31:0] operation_274_2071;
wire signed [31:0] operation_274_2070;
wire signed [31:0] operation_274_2069;
wire signed [31:0] operation_274_2068;
wire signed [31:0] operation_274_2067;
wire signed [31:0] operation_274_2066;
wire signed [31:0] operation_274_2065;
wire signed [31:0] operation_274_2064;
wire signed [31:0] operation_274_2063;
wire signed [31:0] operation_274_2062;
wire signed [31:0] operation_274_2061;
wire signed [31:0] operation_274_2060;
wire signed [31:0] operation_274_2010;
wire signed [31:0] operation_274_2009;
wire signed [31:0] operation_274_1988;
wire signed [31:0] operation_274_1987;
reg [7:0] operation_274_2104_latch;
wire [7:0] operation_274_2104;
reg [7:0] operation_274_2103_latch;
wire [7:0] operation_274_2103;
reg [7:0] operation_274_2102_latch;
wire [7:0] operation_274_2102;
reg [7:0] operation_274_2101_latch;
wire [7:0] operation_274_2101;
reg [7:0] operation_274_2100_latch;
wire [7:0] operation_274_2100;
reg [7:0] operation_274_2099_latch;
wire [7:0] operation_274_2099;
reg [7:0] operation_274_2098_latch;
wire [7:0] operation_274_2098;
reg [7:0] operation_274_2097_latch;
wire [7:0] operation_274_2097;
reg [7:0] operation_274_2096_latch;
wire [7:0] operation_274_2096;
reg [7:0] operation_274_2095_latch;
wire [7:0] operation_274_2095;
reg [7:0] operation_274_2094_latch;
wire [7:0] operation_274_2094;
reg [7:0] operation_274_2093_latch;
wire [7:0] operation_274_2093;
reg [7:0] operation_274_2092_latch;
wire [7:0] operation_274_2092;
reg [7:0] operation_274_2091_latch;
wire [7:0] operation_274_2091;
reg [7:0] operation_274_2090_latch;
wire [7:0] operation_274_2090;
reg [7:0] operation_274_2089_latch;
wire [7:0] operation_274_2089;
wire [7:0] operation_274_2035;
wire [7:0] operation_274_2034;
wire [7:0] operation_274_2033;
wire [7:0] operation_274_2012;
wire [7:0] operation_274_119;
wire [7:0] operation_274_103;
wire [7:0] operation_274_87;
wire [7:0] operation_274_71;
wire [7:0] operation_274_55;
wire [7:0] operation_274_39;
wire [7:0] operation_274_23;
wire [7:0] operation_274_7;
wire [7:0] operation_274_15;
wire [7:0] operation_274_31;
wire [7:0] operation_274_47;
wire [7:0] operation_274_63;
wire [7:0] operation_274_79;
wire [7:0] operation_274_95;
wire [7:0] operation_274_111;
wire [7:0] operation_274_127;
reg signed [31:0] operation_274_2056;
reg signed [31:0] operation_274_2055;
reg signed [31:0] operation_274_2054;
reg signed [31:0] operation_274_2037;
reg signed [31:0] operation_274_118;
reg signed [31:0] operation_274_102;
reg signed [31:0] operation_274_86;
reg signed [31:0] operation_274_70;
reg signed [31:0] operation_274_54;
reg signed [31:0] operation_274_38;
reg signed [31:0] operation_274_22;
reg signed [31:0] operation_274_6;
reg signed [31:0] operation_274_14;
reg signed [31:0] operation_274_30;
reg signed [31:0] operation_274_46;
reg signed [31:0] operation_274_62;
reg signed [31:0] operation_274_78;
reg signed [31:0] operation_274_94;
reg signed [31:0] operation_274_110;
reg signed [31:0] operation_274_126;
wire signed [31:0] operation_274_2078;
wire signed [31:0] operation_274_2077;
wire signed [31:0] operation_274_2076;
wire signed [31:0] operation_274_2059;
wire signed [31:0] operation_274_117;
wire signed [31:0] operation_274_115;
wire signed [31:0] operation_274_101;
wire signed [31:0] operation_274_99;
wire signed [31:0] operation_274_85;
wire signed [31:0] operation_274_83;
wire signed [31:0] operation_274_69;
wire signed [31:0] operation_274_67;
wire signed [31:0] operation_274_53;
wire signed [31:0] operation_274_51;
wire signed [31:0] operation_274_37;
wire signed [31:0] operation_274_35;
wire signed [31:0] operation_274_21;
wire signed [31:0] operation_274_19;
wire signed [31:0] operation_274_5;
wire signed [31:0] operation_274_3;
wire signed [31:0] operation_274_11;
wire signed [31:0] operation_274_13;
wire signed [31:0] operation_274_27;
wire signed [31:0] operation_274_29;
wire signed [31:0] operation_274_43;
wire signed [31:0] operation_274_45;
wire signed [31:0] operation_274_59;
wire signed [31:0] operation_274_61;
wire signed [31:0] operation_274_75;
wire signed [31:0] operation_274_77;
wire signed [31:0] operation_274_91;
wire signed [31:0] operation_274_93;
wire signed [31:0] operation_274_107;
wire signed [31:0] operation_274_109;
wire signed [31:0] operation_274_123;
wire signed [31:0] operation_274_125;
reg [7:0] operation_274_2106_latch;
wire [7:0] operation_274_2106;
reg [7:0] operation_274_2105_latch;
wire [7:0] operation_274_2105;
reg [7:0] operation_274_2088_latch;
wire [7:0] operation_274_2088;
reg [7:0] operation_274_2087_latch;
wire [7:0] operation_274_2087;
wire signed [31:0] operation_274_5601;
wire signed [31:0] operation_274_5597;
wire signed [31:0] operation_274_5592;
wire signed [31:0] operation_274_5587;
wire signed [31:0] operation_274_5582;
wire signed [31:0] operation_274_5577;
wire signed [31:0] operation_274_5572;
wire signed [31:0] operation_274_5567;
wire signed [31:0] operation_274_5562;
wire signed [31:0] operation_274_5557;
wire signed [31:0] operation_274_2119;
wire [127:0] operation_274_124;
wire [127:0] operation_274_122;
reg control_274_follow;
wire control_274_end;
wire control_274_0;
reg control_274_start;
reg control_274_84;
reg control_274_83;
reg control_274_82;
reg control_274_81;
reg control_274_80;
reg control_274_79;
reg control_274_78;
reg control_274_77;
reg control_274_76;
reg control_274_75;
reg control_274_74;
reg control_274_73;
reg control_274_72;
reg control_274_71;
reg control_274_70;
reg control_274_69;
reg control_274_68;
reg control_274_67;
reg control_274_66;
reg control_274_65;
reg control_274_64;
reg control_274_63;
reg control_274_62;
reg control_274_61;
reg control_274_60;
reg control_274_59;
reg control_274_58;
reg control_274_57;
reg control_274_56;
reg control_274_55;
reg control_274_54;
reg control_274_53;
reg control_274_52;
reg control_274_51;
reg control_274_50;
reg control_274_49;
reg control_274_48;
reg control_274_47;
reg control_274_46;
reg control_274_45;
reg control_274_44;
reg control_274_43;
reg control_274_42;
reg control_274_41;
reg control_274_40;
reg control_274_39;
reg control_274_38;
reg control_274_37;
reg control_274_36;
reg control_274_35;
reg control_274_34;
reg control_274_33;
reg control_274_32;
reg control_274_31;
reg control_274_30;
reg control_274_29;
reg control_274_28;
reg control_274_27;
reg control_274_26;
reg control_274_25;
reg control_274_24;
reg control_274_23;
reg control_274_22;
reg control_274_21;
reg control_274_20;
reg control_274_19;
reg control_274_18;
reg control_274_17;
reg control_274_16;
reg control_274_15;
reg control_274_14;
reg control_274_13;
reg control_274_12;
reg control_274_11;
reg control_274_10;
reg control_274_9;
reg control_274_8;
reg control_274_7;
reg control_274_6;
reg control_274_5;
reg control_274_4;
reg control_274_3;
reg control_274_2;
reg control_274_1;
reg [127:0] input_key_274_follow;
wire [127:0] input_key_274;
reg [127:0] input_in_274_follow;
wire [127:0] input_in_274;
reg [7:0] lookup_sbox_0_output;
reg [7:0] sbox_0[256];
wire lookup_sbox_0_enable;
wire [255:0] lookup_sbox_0_0;
reg [7:0] lookup_sbox_1_output;
reg [7:0] sbox_1[256];
wire lookup_sbox_1_enable;
wire [255:0] lookup_sbox_1_0;
reg [7:0] lookup_sbox_2_output;
reg [7:0] sbox_2[256];
wire lookup_sbox_2_enable;
wire [255:0] lookup_sbox_2_0;
reg [7:0] lookup_sbox_3_output;
reg [7:0] sbox_3[256];
wire lookup_sbox_3_enable;
wire [255:0] lookup_sbox_3_0;
reg [7:0] lookup_sbox_4_output;
reg [7:0] sbox_4[256];
wire lookup_sbox_4_enable;
wire [255:0] lookup_sbox_4_0;
reg [7:0] lookup_sbox_5_output;
reg [7:0] sbox_5[256];
wire lookup_sbox_5_enable;
wire [255:0] lookup_sbox_5_0;
reg [7:0] lookup_sbox_6_output;
reg [7:0] sbox_6[256];
wire lookup_sbox_6_enable;
wire [255:0] lookup_sbox_6_0;
reg [7:0] lookup_sbox_7_output;
reg [7:0] sbox_7[256];
wire lookup_sbox_7_enable;
wire [255:0] lookup_sbox_7_0;
reg [7:0] lookup_sbox_8_output;
reg [7:0] sbox_8[256];
wire lookup_sbox_8_enable;
wire [255:0] lookup_sbox_8_0;
reg [7:0] lookup_sbox_9_output;
reg [7:0] sbox_9[256];
wire lookup_sbox_9_enable;
wire [255:0] lookup_sbox_9_0;
reg [7:0] lookup_sbox_10_output;
reg [7:0] sbox_10[256];
wire lookup_sbox_10_enable;
wire [255:0] lookup_sbox_10_0;
reg [7:0] lookup_sbox_11_output;
reg [7:0] sbox_11[256];
wire lookup_sbox_11_enable;
wire [255:0] lookup_sbox_11_0;
reg [7:0] lookup_sbox_12_output;
reg [7:0] sbox_12[256];
wire lookup_sbox_12_enable;
wire [255:0] lookup_sbox_12_0;
reg [7:0] lookup_sbox_13_output;
reg [7:0] sbox_13[256];
wire lookup_sbox_13_enable;
wire [255:0] lookup_sbox_13_0;
reg [7:0] lookup_sbox_14_output;
reg [7:0] sbox_14[256];
wire lookup_sbox_14_enable;
wire [255:0] lookup_sbox_14_0;
reg [7:0] lookup_sbox_15_output;
reg [7:0] sbox_15[256];
wire lookup_sbox_15_enable;
wire [255:0] lookup_sbox_15_0;
reg startfollow;
initial begin
    
    sbox_0[0] = 8'd99;
    sbox_0[1] = 8'd124;
    sbox_0[2] = 8'd119;
    sbox_0[3] = 8'd123;
    sbox_0[4] = 8'd242;
    sbox_0[5] = 8'd107;
    sbox_0[6] = 8'd111;
    sbox_0[7] = 8'd197;
    sbox_0[8] = 8'd48;
    sbox_0[9] = 8'd1;
    sbox_0[10] = 8'd103;
    sbox_0[11] = 8'd43;
    sbox_0[12] = 8'd254;
    sbox_0[13] = 8'd215;
    sbox_0[14] = 8'd171;
    sbox_0[15] = 8'd118;
    sbox_0[16] = 8'd202;
    sbox_0[17] = 8'd130;
    sbox_0[18] = 8'd201;
    sbox_0[19] = 8'd125;
    sbox_0[20] = 8'd250;
    sbox_0[21] = 8'd89;
    sbox_0[22] = 8'd71;
    sbox_0[23] = 8'd240;
    sbox_0[24] = 8'd173;
    sbox_0[25] = 8'd212;
    sbox_0[26] = 8'd162;
    sbox_0[27] = 8'd175;
    sbox_0[28] = 8'd156;
    sbox_0[29] = 8'd164;
    sbox_0[30] = 8'd114;
    sbox_0[31] = 8'd192;
    sbox_0[32] = 8'd183;
    sbox_0[33] = 8'd253;
    sbox_0[34] = 8'd147;
    sbox_0[35] = 8'd38;
    sbox_0[36] = 8'd54;
    sbox_0[37] = 8'd63;
    sbox_0[38] = 8'd247;
    sbox_0[39] = 8'd204;
    sbox_0[40] = 8'd52;
    sbox_0[41] = 8'd165;
    sbox_0[42] = 8'd229;
    sbox_0[43] = 8'd241;
    sbox_0[44] = 8'd113;
    sbox_0[45] = 8'd216;
    sbox_0[46] = 8'd49;
    sbox_0[47] = 8'd21;
    sbox_0[48] = 8'd4;
    sbox_0[49] = 8'd199;
    sbox_0[50] = 8'd35;
    sbox_0[51] = 8'd195;
    sbox_0[52] = 8'd24;
    sbox_0[53] = 8'd150;
    sbox_0[54] = 8'd5;
    sbox_0[55] = 8'd154;
    sbox_0[56] = 8'd7;
    sbox_0[57] = 8'd18;
    sbox_0[58] = 8'd128;
    sbox_0[59] = 8'd226;
    sbox_0[60] = 8'd235;
    sbox_0[61] = 8'd39;
    sbox_0[62] = 8'd178;
    sbox_0[63] = 8'd117;
    sbox_0[64] = 8'd9;
    sbox_0[65] = 8'd131;
    sbox_0[66] = 8'd44;
    sbox_0[67] = 8'd26;
    sbox_0[68] = 8'd27;
    sbox_0[69] = 8'd110;
    sbox_0[70] = 8'd90;
    sbox_0[71] = 8'd160;
    sbox_0[72] = 8'd82;
    sbox_0[73] = 8'd59;
    sbox_0[74] = 8'd214;
    sbox_0[75] = 8'd179;
    sbox_0[76] = 8'd41;
    sbox_0[77] = 8'd227;
    sbox_0[78] = 8'd47;
    sbox_0[79] = 8'd132;
    sbox_0[80] = 8'd83;
    sbox_0[81] = 8'd209;
    sbox_0[82] = 8'd0;
    sbox_0[83] = 8'd237;
    sbox_0[84] = 8'd32;
    sbox_0[85] = 8'd252;
    sbox_0[86] = 8'd177;
    sbox_0[87] = 8'd91;
    sbox_0[88] = 8'd106;
    sbox_0[89] = 8'd203;
    sbox_0[90] = 8'd190;
    sbox_0[91] = 8'd57;
    sbox_0[92] = 8'd74;
    sbox_0[93] = 8'd76;
    sbox_0[94] = 8'd88;
    sbox_0[95] = 8'd207;
    sbox_0[96] = 8'd208;
    sbox_0[97] = 8'd239;
    sbox_0[98] = 8'd170;
    sbox_0[99] = 8'd251;
    sbox_0[100] = 8'd67;
    sbox_0[101] = 8'd77;
    sbox_0[102] = 8'd51;
    sbox_0[103] = 8'd133;
    sbox_0[104] = 8'd69;
    sbox_0[105] = 8'd249;
    sbox_0[106] = 8'd2;
    sbox_0[107] = 8'd127;
    sbox_0[108] = 8'd80;
    sbox_0[109] = 8'd60;
    sbox_0[110] = 8'd159;
    sbox_0[111] = 8'd168;
    sbox_0[112] = 8'd81;
    sbox_0[113] = 8'd163;
    sbox_0[114] = 8'd64;
    sbox_0[115] = 8'd143;
    sbox_0[116] = 8'd146;
    sbox_0[117] = 8'd157;
    sbox_0[118] = 8'd56;
    sbox_0[119] = 8'd245;
    sbox_0[120] = 8'd188;
    sbox_0[121] = 8'd182;
    sbox_0[122] = 8'd218;
    sbox_0[123] = 8'd33;
    sbox_0[124] = 8'd16;
    sbox_0[125] = 8'd255;
    sbox_0[126] = 8'd243;
    sbox_0[127] = 8'd210;
    sbox_0[128] = 8'd205;
    sbox_0[129] = 8'd12;
    sbox_0[130] = 8'd19;
    sbox_0[131] = 8'd236;
    sbox_0[132] = 8'd95;
    sbox_0[133] = 8'd151;
    sbox_0[134] = 8'd68;
    sbox_0[135] = 8'd23;
    sbox_0[136] = 8'd196;
    sbox_0[137] = 8'd167;
    sbox_0[138] = 8'd126;
    sbox_0[139] = 8'd61;
    sbox_0[140] = 8'd100;
    sbox_0[141] = 8'd93;
    sbox_0[142] = 8'd25;
    sbox_0[143] = 8'd115;
    sbox_0[144] = 8'd96;
    sbox_0[145] = 8'd129;
    sbox_0[146] = 8'd79;
    sbox_0[147] = 8'd220;
    sbox_0[148] = 8'd34;
    sbox_0[149] = 8'd42;
    sbox_0[150] = 8'd144;
    sbox_0[151] = 8'd136;
    sbox_0[152] = 8'd70;
    sbox_0[153] = 8'd238;
    sbox_0[154] = 8'd184;
    sbox_0[155] = 8'd20;
    sbox_0[156] = 8'd222;
    sbox_0[157] = 8'd94;
    sbox_0[158] = 8'd11;
    sbox_0[159] = 8'd219;
    sbox_0[160] = 8'd224;
    sbox_0[161] = 8'd50;
    sbox_0[162] = 8'd58;
    sbox_0[163] = 8'd10;
    sbox_0[164] = 8'd73;
    sbox_0[165] = 8'd6;
    sbox_0[166] = 8'd36;
    sbox_0[167] = 8'd92;
    sbox_0[168] = 8'd194;
    sbox_0[169] = 8'd211;
    sbox_0[170] = 8'd172;
    sbox_0[171] = 8'd98;
    sbox_0[172] = 8'd145;
    sbox_0[173] = 8'd149;
    sbox_0[174] = 8'd228;
    sbox_0[175] = 8'd121;
    sbox_0[176] = 8'd231;
    sbox_0[177] = 8'd200;
    sbox_0[178] = 8'd55;
    sbox_0[179] = 8'd109;
    sbox_0[180] = 8'd141;
    sbox_0[181] = 8'd213;
    sbox_0[182] = 8'd78;
    sbox_0[183] = 8'd169;
    sbox_0[184] = 8'd108;
    sbox_0[185] = 8'd86;
    sbox_0[186] = 8'd244;
    sbox_0[187] = 8'd234;
    sbox_0[188] = 8'd101;
    sbox_0[189] = 8'd122;
    sbox_0[190] = 8'd174;
    sbox_0[191] = 8'd8;
    sbox_0[192] = 8'd186;
    sbox_0[193] = 8'd120;
    sbox_0[194] = 8'd37;
    sbox_0[195] = 8'd46;
    sbox_0[196] = 8'd28;
    sbox_0[197] = 8'd166;
    sbox_0[198] = 8'd180;
    sbox_0[199] = 8'd198;
    sbox_0[200] = 8'd232;
    sbox_0[201] = 8'd221;
    sbox_0[202] = 8'd116;
    sbox_0[203] = 8'd31;
    sbox_0[204] = 8'd75;
    sbox_0[205] = 8'd189;
    sbox_0[206] = 8'd139;
    sbox_0[207] = 8'd138;
    sbox_0[208] = 8'd112;
    sbox_0[209] = 8'd62;
    sbox_0[210] = 8'd181;
    sbox_0[211] = 8'd102;
    sbox_0[212] = 8'd72;
    sbox_0[213] = 8'd3;
    sbox_0[214] = 8'd246;
    sbox_0[215] = 8'd14;
    sbox_0[216] = 8'd97;
    sbox_0[217] = 8'd53;
    sbox_0[218] = 8'd87;
    sbox_0[219] = 8'd185;
    sbox_0[220] = 8'd134;
    sbox_0[221] = 8'd193;
    sbox_0[222] = 8'd29;
    sbox_0[223] = 8'd158;
    sbox_0[224] = 8'd225;
    sbox_0[225] = 8'd248;
    sbox_0[226] = 8'd152;
    sbox_0[227] = 8'd17;
    sbox_0[228] = 8'd105;
    sbox_0[229] = 8'd217;
    sbox_0[230] = 8'd142;
    sbox_0[231] = 8'd148;
    sbox_0[232] = 8'd155;
    sbox_0[233] = 8'd30;
    sbox_0[234] = 8'd135;
    sbox_0[235] = 8'd233;
    sbox_0[236] = 8'd206;
    sbox_0[237] = 8'd85;
    sbox_0[238] = 8'd40;
    sbox_0[239] = 8'd223;
    sbox_0[240] = 8'd140;
    sbox_0[241] = 8'd161;
    sbox_0[242] = 8'd137;
    sbox_0[243] = 8'd13;
    sbox_0[244] = 8'd191;
    sbox_0[245] = 8'd230;
    sbox_0[246] = 8'd66;
    sbox_0[247] = 8'd104;
    sbox_0[248] = 8'd65;
    sbox_0[249] = 8'd153;
    sbox_0[250] = 8'd45;
    sbox_0[251] = 8'd15;
    sbox_0[252] = 8'd176;
    sbox_0[253] = 8'd84;
    sbox_0[254] = 8'd187;
    sbox_0[255] = 8'd22;
    sbox_1[0] = 8'd99;
    sbox_1[1] = 8'd124;
    sbox_1[2] = 8'd119;
    sbox_1[3] = 8'd123;
    sbox_1[4] = 8'd242;
    sbox_1[5] = 8'd107;
    sbox_1[6] = 8'd111;
    sbox_1[7] = 8'd197;
    sbox_1[8] = 8'd48;
    sbox_1[9] = 8'd1;
    sbox_1[10] = 8'd103;
    sbox_1[11] = 8'd43;
    sbox_1[12] = 8'd254;
    sbox_1[13] = 8'd215;
    sbox_1[14] = 8'd171;
    sbox_1[15] = 8'd118;
    sbox_1[16] = 8'd202;
    sbox_1[17] = 8'd130;
    sbox_1[18] = 8'd201;
    sbox_1[19] = 8'd125;
    sbox_1[20] = 8'd250;
    sbox_1[21] = 8'd89;
    sbox_1[22] = 8'd71;
    sbox_1[23] = 8'd240;
    sbox_1[24] = 8'd173;
    sbox_1[25] = 8'd212;
    sbox_1[26] = 8'd162;
    sbox_1[27] = 8'd175;
    sbox_1[28] = 8'd156;
    sbox_1[29] = 8'd164;
    sbox_1[30] = 8'd114;
    sbox_1[31] = 8'd192;
    sbox_1[32] = 8'd183;
    sbox_1[33] = 8'd253;
    sbox_1[34] = 8'd147;
    sbox_1[35] = 8'd38;
    sbox_1[36] = 8'd54;
    sbox_1[37] = 8'd63;
    sbox_1[38] = 8'd247;
    sbox_1[39] = 8'd204;
    sbox_1[40] = 8'd52;
    sbox_1[41] = 8'd165;
    sbox_1[42] = 8'd229;
    sbox_1[43] = 8'd241;
    sbox_1[44] = 8'd113;
    sbox_1[45] = 8'd216;
    sbox_1[46] = 8'd49;
    sbox_1[47] = 8'd21;
    sbox_1[48] = 8'd4;
    sbox_1[49] = 8'd199;
    sbox_1[50] = 8'd35;
    sbox_1[51] = 8'd195;
    sbox_1[52] = 8'd24;
    sbox_1[53] = 8'd150;
    sbox_1[54] = 8'd5;
    sbox_1[55] = 8'd154;
    sbox_1[56] = 8'd7;
    sbox_1[57] = 8'd18;
    sbox_1[58] = 8'd128;
    sbox_1[59] = 8'd226;
    sbox_1[60] = 8'd235;
    sbox_1[61] = 8'd39;
    sbox_1[62] = 8'd178;
    sbox_1[63] = 8'd117;
    sbox_1[64] = 8'd9;
    sbox_1[65] = 8'd131;
    sbox_1[66] = 8'd44;
    sbox_1[67] = 8'd26;
    sbox_1[68] = 8'd27;
    sbox_1[69] = 8'd110;
    sbox_1[70] = 8'd90;
    sbox_1[71] = 8'd160;
    sbox_1[72] = 8'd82;
    sbox_1[73] = 8'd59;
    sbox_1[74] = 8'd214;
    sbox_1[75] = 8'd179;
    sbox_1[76] = 8'd41;
    sbox_1[77] = 8'd227;
    sbox_1[78] = 8'd47;
    sbox_1[79] = 8'd132;
    sbox_1[80] = 8'd83;
    sbox_1[81] = 8'd209;
    sbox_1[82] = 8'd0;
    sbox_1[83] = 8'd237;
    sbox_1[84] = 8'd32;
    sbox_1[85] = 8'd252;
    sbox_1[86] = 8'd177;
    sbox_1[87] = 8'd91;
    sbox_1[88] = 8'd106;
    sbox_1[89] = 8'd203;
    sbox_1[90] = 8'd190;
    sbox_1[91] = 8'd57;
    sbox_1[92] = 8'd74;
    sbox_1[93] = 8'd76;
    sbox_1[94] = 8'd88;
    sbox_1[95] = 8'd207;
    sbox_1[96] = 8'd208;
    sbox_1[97] = 8'd239;
    sbox_1[98] = 8'd170;
    sbox_1[99] = 8'd251;
    sbox_1[100] = 8'd67;
    sbox_1[101] = 8'd77;
    sbox_1[102] = 8'd51;
    sbox_1[103] = 8'd133;
    sbox_1[104] = 8'd69;
    sbox_1[105] = 8'd249;
    sbox_1[106] = 8'd2;
    sbox_1[107] = 8'd127;
    sbox_1[108] = 8'd80;
    sbox_1[109] = 8'd60;
    sbox_1[110] = 8'd159;
    sbox_1[111] = 8'd168;
    sbox_1[112] = 8'd81;
    sbox_1[113] = 8'd163;
    sbox_1[114] = 8'd64;
    sbox_1[115] = 8'd143;
    sbox_1[116] = 8'd146;
    sbox_1[117] = 8'd157;
    sbox_1[118] = 8'd56;
    sbox_1[119] = 8'd245;
    sbox_1[120] = 8'd188;
    sbox_1[121] = 8'd182;
    sbox_1[122] = 8'd218;
    sbox_1[123] = 8'd33;
    sbox_1[124] = 8'd16;
    sbox_1[125] = 8'd255;
    sbox_1[126] = 8'd243;
    sbox_1[127] = 8'd210;
    sbox_1[128] = 8'd205;
    sbox_1[129] = 8'd12;
    sbox_1[130] = 8'd19;
    sbox_1[131] = 8'd236;
    sbox_1[132] = 8'd95;
    sbox_1[133] = 8'd151;
    sbox_1[134] = 8'd68;
    sbox_1[135] = 8'd23;
    sbox_1[136] = 8'd196;
    sbox_1[137] = 8'd167;
    sbox_1[138] = 8'd126;
    sbox_1[139] = 8'd61;
    sbox_1[140] = 8'd100;
    sbox_1[141] = 8'd93;
    sbox_1[142] = 8'd25;
    sbox_1[143] = 8'd115;
    sbox_1[144] = 8'd96;
    sbox_1[145] = 8'd129;
    sbox_1[146] = 8'd79;
    sbox_1[147] = 8'd220;
    sbox_1[148] = 8'd34;
    sbox_1[149] = 8'd42;
    sbox_1[150] = 8'd144;
    sbox_1[151] = 8'd136;
    sbox_1[152] = 8'd70;
    sbox_1[153] = 8'd238;
    sbox_1[154] = 8'd184;
    sbox_1[155] = 8'd20;
    sbox_1[156] = 8'd222;
    sbox_1[157] = 8'd94;
    sbox_1[158] = 8'd11;
    sbox_1[159] = 8'd219;
    sbox_1[160] = 8'd224;
    sbox_1[161] = 8'd50;
    sbox_1[162] = 8'd58;
    sbox_1[163] = 8'd10;
    sbox_1[164] = 8'd73;
    sbox_1[165] = 8'd6;
    sbox_1[166] = 8'd36;
    sbox_1[167] = 8'd92;
    sbox_1[168] = 8'd194;
    sbox_1[169] = 8'd211;
    sbox_1[170] = 8'd172;
    sbox_1[171] = 8'd98;
    sbox_1[172] = 8'd145;
    sbox_1[173] = 8'd149;
    sbox_1[174] = 8'd228;
    sbox_1[175] = 8'd121;
    sbox_1[176] = 8'd231;
    sbox_1[177] = 8'd200;
    sbox_1[178] = 8'd55;
    sbox_1[179] = 8'd109;
    sbox_1[180] = 8'd141;
    sbox_1[181] = 8'd213;
    sbox_1[182] = 8'd78;
    sbox_1[183] = 8'd169;
    sbox_1[184] = 8'd108;
    sbox_1[185] = 8'd86;
    sbox_1[186] = 8'd244;
    sbox_1[187] = 8'd234;
    sbox_1[188] = 8'd101;
    sbox_1[189] = 8'd122;
    sbox_1[190] = 8'd174;
    sbox_1[191] = 8'd8;
    sbox_1[192] = 8'd186;
    sbox_1[193] = 8'd120;
    sbox_1[194] = 8'd37;
    sbox_1[195] = 8'd46;
    sbox_1[196] = 8'd28;
    sbox_1[197] = 8'd166;
    sbox_1[198] = 8'd180;
    sbox_1[199] = 8'd198;
    sbox_1[200] = 8'd232;
    sbox_1[201] = 8'd221;
    sbox_1[202] = 8'd116;
    sbox_1[203] = 8'd31;
    sbox_1[204] = 8'd75;
    sbox_1[205] = 8'd189;
    sbox_1[206] = 8'd139;
    sbox_1[207] = 8'd138;
    sbox_1[208] = 8'd112;
    sbox_1[209] = 8'd62;
    sbox_1[210] = 8'd181;
    sbox_1[211] = 8'd102;
    sbox_1[212] = 8'd72;
    sbox_1[213] = 8'd3;
    sbox_1[214] = 8'd246;
    sbox_1[215] = 8'd14;
    sbox_1[216] = 8'd97;
    sbox_1[217] = 8'd53;
    sbox_1[218] = 8'd87;
    sbox_1[219] = 8'd185;
    sbox_1[220] = 8'd134;
    sbox_1[221] = 8'd193;
    sbox_1[222] = 8'd29;
    sbox_1[223] = 8'd158;
    sbox_1[224] = 8'd225;
    sbox_1[225] = 8'd248;
    sbox_1[226] = 8'd152;
    sbox_1[227] = 8'd17;
    sbox_1[228] = 8'd105;
    sbox_1[229] = 8'd217;
    sbox_1[230] = 8'd142;
    sbox_1[231] = 8'd148;
    sbox_1[232] = 8'd155;
    sbox_1[233] = 8'd30;
    sbox_1[234] = 8'd135;
    sbox_1[235] = 8'd233;
    sbox_1[236] = 8'd206;
    sbox_1[237] = 8'd85;
    sbox_1[238] = 8'd40;
    sbox_1[239] = 8'd223;
    sbox_1[240] = 8'd140;
    sbox_1[241] = 8'd161;
    sbox_1[242] = 8'd137;
    sbox_1[243] = 8'd13;
    sbox_1[244] = 8'd191;
    sbox_1[245] = 8'd230;
    sbox_1[246] = 8'd66;
    sbox_1[247] = 8'd104;
    sbox_1[248] = 8'd65;
    sbox_1[249] = 8'd153;
    sbox_1[250] = 8'd45;
    sbox_1[251] = 8'd15;
    sbox_1[252] = 8'd176;
    sbox_1[253] = 8'd84;
    sbox_1[254] = 8'd187;
    sbox_1[255] = 8'd22;
    sbox_2[0] = 8'd99;
    sbox_2[1] = 8'd124;
    sbox_2[2] = 8'd119;
    sbox_2[3] = 8'd123;
    sbox_2[4] = 8'd242;
    sbox_2[5] = 8'd107;
    sbox_2[6] = 8'd111;
    sbox_2[7] = 8'd197;
    sbox_2[8] = 8'd48;
    sbox_2[9] = 8'd1;
    sbox_2[10] = 8'd103;
    sbox_2[11] = 8'd43;
    sbox_2[12] = 8'd254;
    sbox_2[13] = 8'd215;
    sbox_2[14] = 8'd171;
    sbox_2[15] = 8'd118;
    sbox_2[16] = 8'd202;
    sbox_2[17] = 8'd130;
    sbox_2[18] = 8'd201;
    sbox_2[19] = 8'd125;
    sbox_2[20] = 8'd250;
    sbox_2[21] = 8'd89;
    sbox_2[22] = 8'd71;
    sbox_2[23] = 8'd240;
    sbox_2[24] = 8'd173;
    sbox_2[25] = 8'd212;
    sbox_2[26] = 8'd162;
    sbox_2[27] = 8'd175;
    sbox_2[28] = 8'd156;
    sbox_2[29] = 8'd164;
    sbox_2[30] = 8'd114;
    sbox_2[31] = 8'd192;
    sbox_2[32] = 8'd183;
    sbox_2[33] = 8'd253;
    sbox_2[34] = 8'd147;
    sbox_2[35] = 8'd38;
    sbox_2[36] = 8'd54;
    sbox_2[37] = 8'd63;
    sbox_2[38] = 8'd247;
    sbox_2[39] = 8'd204;
    sbox_2[40] = 8'd52;
    sbox_2[41] = 8'd165;
    sbox_2[42] = 8'd229;
    sbox_2[43] = 8'd241;
    sbox_2[44] = 8'd113;
    sbox_2[45] = 8'd216;
    sbox_2[46] = 8'd49;
    sbox_2[47] = 8'd21;
    sbox_2[48] = 8'd4;
    sbox_2[49] = 8'd199;
    sbox_2[50] = 8'd35;
    sbox_2[51] = 8'd195;
    sbox_2[52] = 8'd24;
    sbox_2[53] = 8'd150;
    sbox_2[54] = 8'd5;
    sbox_2[55] = 8'd154;
    sbox_2[56] = 8'd7;
    sbox_2[57] = 8'd18;
    sbox_2[58] = 8'd128;
    sbox_2[59] = 8'd226;
    sbox_2[60] = 8'd235;
    sbox_2[61] = 8'd39;
    sbox_2[62] = 8'd178;
    sbox_2[63] = 8'd117;
    sbox_2[64] = 8'd9;
    sbox_2[65] = 8'd131;
    sbox_2[66] = 8'd44;
    sbox_2[67] = 8'd26;
    sbox_2[68] = 8'd27;
    sbox_2[69] = 8'd110;
    sbox_2[70] = 8'd90;
    sbox_2[71] = 8'd160;
    sbox_2[72] = 8'd82;
    sbox_2[73] = 8'd59;
    sbox_2[74] = 8'd214;
    sbox_2[75] = 8'd179;
    sbox_2[76] = 8'd41;
    sbox_2[77] = 8'd227;
    sbox_2[78] = 8'd47;
    sbox_2[79] = 8'd132;
    sbox_2[80] = 8'd83;
    sbox_2[81] = 8'd209;
    sbox_2[82] = 8'd0;
    sbox_2[83] = 8'd237;
    sbox_2[84] = 8'd32;
    sbox_2[85] = 8'd252;
    sbox_2[86] = 8'd177;
    sbox_2[87] = 8'd91;
    sbox_2[88] = 8'd106;
    sbox_2[89] = 8'd203;
    sbox_2[90] = 8'd190;
    sbox_2[91] = 8'd57;
    sbox_2[92] = 8'd74;
    sbox_2[93] = 8'd76;
    sbox_2[94] = 8'd88;
    sbox_2[95] = 8'd207;
    sbox_2[96] = 8'd208;
    sbox_2[97] = 8'd239;
    sbox_2[98] = 8'd170;
    sbox_2[99] = 8'd251;
    sbox_2[100] = 8'd67;
    sbox_2[101] = 8'd77;
    sbox_2[102] = 8'd51;
    sbox_2[103] = 8'd133;
    sbox_2[104] = 8'd69;
    sbox_2[105] = 8'd249;
    sbox_2[106] = 8'd2;
    sbox_2[107] = 8'd127;
    sbox_2[108] = 8'd80;
    sbox_2[109] = 8'd60;
    sbox_2[110] = 8'd159;
    sbox_2[111] = 8'd168;
    sbox_2[112] = 8'd81;
    sbox_2[113] = 8'd163;
    sbox_2[114] = 8'd64;
    sbox_2[115] = 8'd143;
    sbox_2[116] = 8'd146;
    sbox_2[117] = 8'd157;
    sbox_2[118] = 8'd56;
    sbox_2[119] = 8'd245;
    sbox_2[120] = 8'd188;
    sbox_2[121] = 8'd182;
    sbox_2[122] = 8'd218;
    sbox_2[123] = 8'd33;
    sbox_2[124] = 8'd16;
    sbox_2[125] = 8'd255;
    sbox_2[126] = 8'd243;
    sbox_2[127] = 8'd210;
    sbox_2[128] = 8'd205;
    sbox_2[129] = 8'd12;
    sbox_2[130] = 8'd19;
    sbox_2[131] = 8'd236;
    sbox_2[132] = 8'd95;
    sbox_2[133] = 8'd151;
    sbox_2[134] = 8'd68;
    sbox_2[135] = 8'd23;
    sbox_2[136] = 8'd196;
    sbox_2[137] = 8'd167;
    sbox_2[138] = 8'd126;
    sbox_2[139] = 8'd61;
    sbox_2[140] = 8'd100;
    sbox_2[141] = 8'd93;
    sbox_2[142] = 8'd25;
    sbox_2[143] = 8'd115;
    sbox_2[144] = 8'd96;
    sbox_2[145] = 8'd129;
    sbox_2[146] = 8'd79;
    sbox_2[147] = 8'd220;
    sbox_2[148] = 8'd34;
    sbox_2[149] = 8'd42;
    sbox_2[150] = 8'd144;
    sbox_2[151] = 8'd136;
    sbox_2[152] = 8'd70;
    sbox_2[153] = 8'd238;
    sbox_2[154] = 8'd184;
    sbox_2[155] = 8'd20;
    sbox_2[156] = 8'd222;
    sbox_2[157] = 8'd94;
    sbox_2[158] = 8'd11;
    sbox_2[159] = 8'd219;
    sbox_2[160] = 8'd224;
    sbox_2[161] = 8'd50;
    sbox_2[162] = 8'd58;
    sbox_2[163] = 8'd10;
    sbox_2[164] = 8'd73;
    sbox_2[165] = 8'd6;
    sbox_2[166] = 8'd36;
    sbox_2[167] = 8'd92;
    sbox_2[168] = 8'd194;
    sbox_2[169] = 8'd211;
    sbox_2[170] = 8'd172;
    sbox_2[171] = 8'd98;
    sbox_2[172] = 8'd145;
    sbox_2[173] = 8'd149;
    sbox_2[174] = 8'd228;
    sbox_2[175] = 8'd121;
    sbox_2[176] = 8'd231;
    sbox_2[177] = 8'd200;
    sbox_2[178] = 8'd55;
    sbox_2[179] = 8'd109;
    sbox_2[180] = 8'd141;
    sbox_2[181] = 8'd213;
    sbox_2[182] = 8'd78;
    sbox_2[183] = 8'd169;
    sbox_2[184] = 8'd108;
    sbox_2[185] = 8'd86;
    sbox_2[186] = 8'd244;
    sbox_2[187] = 8'd234;
    sbox_2[188] = 8'd101;
    sbox_2[189] = 8'd122;
    sbox_2[190] = 8'd174;
    sbox_2[191] = 8'd8;
    sbox_2[192] = 8'd186;
    sbox_2[193] = 8'd120;
    sbox_2[194] = 8'd37;
    sbox_2[195] = 8'd46;
    sbox_2[196] = 8'd28;
    sbox_2[197] = 8'd166;
    sbox_2[198] = 8'd180;
    sbox_2[199] = 8'd198;
    sbox_2[200] = 8'd232;
    sbox_2[201] = 8'd221;
    sbox_2[202] = 8'd116;
    sbox_2[203] = 8'd31;
    sbox_2[204] = 8'd75;
    sbox_2[205] = 8'd189;
    sbox_2[206] = 8'd139;
    sbox_2[207] = 8'd138;
    sbox_2[208] = 8'd112;
    sbox_2[209] = 8'd62;
    sbox_2[210] = 8'd181;
    sbox_2[211] = 8'd102;
    sbox_2[212] = 8'd72;
    sbox_2[213] = 8'd3;
    sbox_2[214] = 8'd246;
    sbox_2[215] = 8'd14;
    sbox_2[216] = 8'd97;
    sbox_2[217] = 8'd53;
    sbox_2[218] = 8'd87;
    sbox_2[219] = 8'd185;
    sbox_2[220] = 8'd134;
    sbox_2[221] = 8'd193;
    sbox_2[222] = 8'd29;
    sbox_2[223] = 8'd158;
    sbox_2[224] = 8'd225;
    sbox_2[225] = 8'd248;
    sbox_2[226] = 8'd152;
    sbox_2[227] = 8'd17;
    sbox_2[228] = 8'd105;
    sbox_2[229] = 8'd217;
    sbox_2[230] = 8'd142;
    sbox_2[231] = 8'd148;
    sbox_2[232] = 8'd155;
    sbox_2[233] = 8'd30;
    sbox_2[234] = 8'd135;
    sbox_2[235] = 8'd233;
    sbox_2[236] = 8'd206;
    sbox_2[237] = 8'd85;
    sbox_2[238] = 8'd40;
    sbox_2[239] = 8'd223;
    sbox_2[240] = 8'd140;
    sbox_2[241] = 8'd161;
    sbox_2[242] = 8'd137;
    sbox_2[243] = 8'd13;
    sbox_2[244] = 8'd191;
    sbox_2[245] = 8'd230;
    sbox_2[246] = 8'd66;
    sbox_2[247] = 8'd104;
    sbox_2[248] = 8'd65;
    sbox_2[249] = 8'd153;
    sbox_2[250] = 8'd45;
    sbox_2[251] = 8'd15;
    sbox_2[252] = 8'd176;
    sbox_2[253] = 8'd84;
    sbox_2[254] = 8'd187;
    sbox_2[255] = 8'd22;
    sbox_3[0] = 8'd99;
    sbox_3[1] = 8'd124;
    sbox_3[2] = 8'd119;
    sbox_3[3] = 8'd123;
    sbox_3[4] = 8'd242;
    sbox_3[5] = 8'd107;
    sbox_3[6] = 8'd111;
    sbox_3[7] = 8'd197;
    sbox_3[8] = 8'd48;
    sbox_3[9] = 8'd1;
    sbox_3[10] = 8'd103;
    sbox_3[11] = 8'd43;
    sbox_3[12] = 8'd254;
    sbox_3[13] = 8'd215;
    sbox_3[14] = 8'd171;
    sbox_3[15] = 8'd118;
    sbox_3[16] = 8'd202;
    sbox_3[17] = 8'd130;
    sbox_3[18] = 8'd201;
    sbox_3[19] = 8'd125;
    sbox_3[20] = 8'd250;
    sbox_3[21] = 8'd89;
    sbox_3[22] = 8'd71;
    sbox_3[23] = 8'd240;
    sbox_3[24] = 8'd173;
    sbox_3[25] = 8'd212;
    sbox_3[26] = 8'd162;
    sbox_3[27] = 8'd175;
    sbox_3[28] = 8'd156;
    sbox_3[29] = 8'd164;
    sbox_3[30] = 8'd114;
    sbox_3[31] = 8'd192;
    sbox_3[32] = 8'd183;
    sbox_3[33] = 8'd253;
    sbox_3[34] = 8'd147;
    sbox_3[35] = 8'd38;
    sbox_3[36] = 8'd54;
    sbox_3[37] = 8'd63;
    sbox_3[38] = 8'd247;
    sbox_3[39] = 8'd204;
    sbox_3[40] = 8'd52;
    sbox_3[41] = 8'd165;
    sbox_3[42] = 8'd229;
    sbox_3[43] = 8'd241;
    sbox_3[44] = 8'd113;
    sbox_3[45] = 8'd216;
    sbox_3[46] = 8'd49;
    sbox_3[47] = 8'd21;
    sbox_3[48] = 8'd4;
    sbox_3[49] = 8'd199;
    sbox_3[50] = 8'd35;
    sbox_3[51] = 8'd195;
    sbox_3[52] = 8'd24;
    sbox_3[53] = 8'd150;
    sbox_3[54] = 8'd5;
    sbox_3[55] = 8'd154;
    sbox_3[56] = 8'd7;
    sbox_3[57] = 8'd18;
    sbox_3[58] = 8'd128;
    sbox_3[59] = 8'd226;
    sbox_3[60] = 8'd235;
    sbox_3[61] = 8'd39;
    sbox_3[62] = 8'd178;
    sbox_3[63] = 8'd117;
    sbox_3[64] = 8'd9;
    sbox_3[65] = 8'd131;
    sbox_3[66] = 8'd44;
    sbox_3[67] = 8'd26;
    sbox_3[68] = 8'd27;
    sbox_3[69] = 8'd110;
    sbox_3[70] = 8'd90;
    sbox_3[71] = 8'd160;
    sbox_3[72] = 8'd82;
    sbox_3[73] = 8'd59;
    sbox_3[74] = 8'd214;
    sbox_3[75] = 8'd179;
    sbox_3[76] = 8'd41;
    sbox_3[77] = 8'd227;
    sbox_3[78] = 8'd47;
    sbox_3[79] = 8'd132;
    sbox_3[80] = 8'd83;
    sbox_3[81] = 8'd209;
    sbox_3[82] = 8'd0;
    sbox_3[83] = 8'd237;
    sbox_3[84] = 8'd32;
    sbox_3[85] = 8'd252;
    sbox_3[86] = 8'd177;
    sbox_3[87] = 8'd91;
    sbox_3[88] = 8'd106;
    sbox_3[89] = 8'd203;
    sbox_3[90] = 8'd190;
    sbox_3[91] = 8'd57;
    sbox_3[92] = 8'd74;
    sbox_3[93] = 8'd76;
    sbox_3[94] = 8'd88;
    sbox_3[95] = 8'd207;
    sbox_3[96] = 8'd208;
    sbox_3[97] = 8'd239;
    sbox_3[98] = 8'd170;
    sbox_3[99] = 8'd251;
    sbox_3[100] = 8'd67;
    sbox_3[101] = 8'd77;
    sbox_3[102] = 8'd51;
    sbox_3[103] = 8'd133;
    sbox_3[104] = 8'd69;
    sbox_3[105] = 8'd249;
    sbox_3[106] = 8'd2;
    sbox_3[107] = 8'd127;
    sbox_3[108] = 8'd80;
    sbox_3[109] = 8'd60;
    sbox_3[110] = 8'd159;
    sbox_3[111] = 8'd168;
    sbox_3[112] = 8'd81;
    sbox_3[113] = 8'd163;
    sbox_3[114] = 8'd64;
    sbox_3[115] = 8'd143;
    sbox_3[116] = 8'd146;
    sbox_3[117] = 8'd157;
    sbox_3[118] = 8'd56;
    sbox_3[119] = 8'd245;
    sbox_3[120] = 8'd188;
    sbox_3[121] = 8'd182;
    sbox_3[122] = 8'd218;
    sbox_3[123] = 8'd33;
    sbox_3[124] = 8'd16;
    sbox_3[125] = 8'd255;
    sbox_3[126] = 8'd243;
    sbox_3[127] = 8'd210;
    sbox_3[128] = 8'd205;
    sbox_3[129] = 8'd12;
    sbox_3[130] = 8'd19;
    sbox_3[131] = 8'd236;
    sbox_3[132] = 8'd95;
    sbox_3[133] = 8'd151;
    sbox_3[134] = 8'd68;
    sbox_3[135] = 8'd23;
    sbox_3[136] = 8'd196;
    sbox_3[137] = 8'd167;
    sbox_3[138] = 8'd126;
    sbox_3[139] = 8'd61;
    sbox_3[140] = 8'd100;
    sbox_3[141] = 8'd93;
    sbox_3[142] = 8'd25;
    sbox_3[143] = 8'd115;
    sbox_3[144] = 8'd96;
    sbox_3[145] = 8'd129;
    sbox_3[146] = 8'd79;
    sbox_3[147] = 8'd220;
    sbox_3[148] = 8'd34;
    sbox_3[149] = 8'd42;
    sbox_3[150] = 8'd144;
    sbox_3[151] = 8'd136;
    sbox_3[152] = 8'd70;
    sbox_3[153] = 8'd238;
    sbox_3[154] = 8'd184;
    sbox_3[155] = 8'd20;
    sbox_3[156] = 8'd222;
    sbox_3[157] = 8'd94;
    sbox_3[158] = 8'd11;
    sbox_3[159] = 8'd219;
    sbox_3[160] = 8'd224;
    sbox_3[161] = 8'd50;
    sbox_3[162] = 8'd58;
    sbox_3[163] = 8'd10;
    sbox_3[164] = 8'd73;
    sbox_3[165] = 8'd6;
    sbox_3[166] = 8'd36;
    sbox_3[167] = 8'd92;
    sbox_3[168] = 8'd194;
    sbox_3[169] = 8'd211;
    sbox_3[170] = 8'd172;
    sbox_3[171] = 8'd98;
    sbox_3[172] = 8'd145;
    sbox_3[173] = 8'd149;
    sbox_3[174] = 8'd228;
    sbox_3[175] = 8'd121;
    sbox_3[176] = 8'd231;
    sbox_3[177] = 8'd200;
    sbox_3[178] = 8'd55;
    sbox_3[179] = 8'd109;
    sbox_3[180] = 8'd141;
    sbox_3[181] = 8'd213;
    sbox_3[182] = 8'd78;
    sbox_3[183] = 8'd169;
    sbox_3[184] = 8'd108;
    sbox_3[185] = 8'd86;
    sbox_3[186] = 8'd244;
    sbox_3[187] = 8'd234;
    sbox_3[188] = 8'd101;
    sbox_3[189] = 8'd122;
    sbox_3[190] = 8'd174;
    sbox_3[191] = 8'd8;
    sbox_3[192] = 8'd186;
    sbox_3[193] = 8'd120;
    sbox_3[194] = 8'd37;
    sbox_3[195] = 8'd46;
    sbox_3[196] = 8'd28;
    sbox_3[197] = 8'd166;
    sbox_3[198] = 8'd180;
    sbox_3[199] = 8'd198;
    sbox_3[200] = 8'd232;
    sbox_3[201] = 8'd221;
    sbox_3[202] = 8'd116;
    sbox_3[203] = 8'd31;
    sbox_3[204] = 8'd75;
    sbox_3[205] = 8'd189;
    sbox_3[206] = 8'd139;
    sbox_3[207] = 8'd138;
    sbox_3[208] = 8'd112;
    sbox_3[209] = 8'd62;
    sbox_3[210] = 8'd181;
    sbox_3[211] = 8'd102;
    sbox_3[212] = 8'd72;
    sbox_3[213] = 8'd3;
    sbox_3[214] = 8'd246;
    sbox_3[215] = 8'd14;
    sbox_3[216] = 8'd97;
    sbox_3[217] = 8'd53;
    sbox_3[218] = 8'd87;
    sbox_3[219] = 8'd185;
    sbox_3[220] = 8'd134;
    sbox_3[221] = 8'd193;
    sbox_3[222] = 8'd29;
    sbox_3[223] = 8'd158;
    sbox_3[224] = 8'd225;
    sbox_3[225] = 8'd248;
    sbox_3[226] = 8'd152;
    sbox_3[227] = 8'd17;
    sbox_3[228] = 8'd105;
    sbox_3[229] = 8'd217;
    sbox_3[230] = 8'd142;
    sbox_3[231] = 8'd148;
    sbox_3[232] = 8'd155;
    sbox_3[233] = 8'd30;
    sbox_3[234] = 8'd135;
    sbox_3[235] = 8'd233;
    sbox_3[236] = 8'd206;
    sbox_3[237] = 8'd85;
    sbox_3[238] = 8'd40;
    sbox_3[239] = 8'd223;
    sbox_3[240] = 8'd140;
    sbox_3[241] = 8'd161;
    sbox_3[242] = 8'd137;
    sbox_3[243] = 8'd13;
    sbox_3[244] = 8'd191;
    sbox_3[245] = 8'd230;
    sbox_3[246] = 8'd66;
    sbox_3[247] = 8'd104;
    sbox_3[248] = 8'd65;
    sbox_3[249] = 8'd153;
    sbox_3[250] = 8'd45;
    sbox_3[251] = 8'd15;
    sbox_3[252] = 8'd176;
    sbox_3[253] = 8'd84;
    sbox_3[254] = 8'd187;
    sbox_3[255] = 8'd22;
    sbox_4[0] = 8'd99;
    sbox_4[1] = 8'd124;
    sbox_4[2] = 8'd119;
    sbox_4[3] = 8'd123;
    sbox_4[4] = 8'd242;
    sbox_4[5] = 8'd107;
    sbox_4[6] = 8'd111;
    sbox_4[7] = 8'd197;
    sbox_4[8] = 8'd48;
    sbox_4[9] = 8'd1;
    sbox_4[10] = 8'd103;
    sbox_4[11] = 8'd43;
    sbox_4[12] = 8'd254;
    sbox_4[13] = 8'd215;
    sbox_4[14] = 8'd171;
    sbox_4[15] = 8'd118;
    sbox_4[16] = 8'd202;
    sbox_4[17] = 8'd130;
    sbox_4[18] = 8'd201;
    sbox_4[19] = 8'd125;
    sbox_4[20] = 8'd250;
    sbox_4[21] = 8'd89;
    sbox_4[22] = 8'd71;
    sbox_4[23] = 8'd240;
    sbox_4[24] = 8'd173;
    sbox_4[25] = 8'd212;
    sbox_4[26] = 8'd162;
    sbox_4[27] = 8'd175;
    sbox_4[28] = 8'd156;
    sbox_4[29] = 8'd164;
    sbox_4[30] = 8'd114;
    sbox_4[31] = 8'd192;
    sbox_4[32] = 8'd183;
    sbox_4[33] = 8'd253;
    sbox_4[34] = 8'd147;
    sbox_4[35] = 8'd38;
    sbox_4[36] = 8'd54;
    sbox_4[37] = 8'd63;
    sbox_4[38] = 8'd247;
    sbox_4[39] = 8'd204;
    sbox_4[40] = 8'd52;
    sbox_4[41] = 8'd165;
    sbox_4[42] = 8'd229;
    sbox_4[43] = 8'd241;
    sbox_4[44] = 8'd113;
    sbox_4[45] = 8'd216;
    sbox_4[46] = 8'd49;
    sbox_4[47] = 8'd21;
    sbox_4[48] = 8'd4;
    sbox_4[49] = 8'd199;
    sbox_4[50] = 8'd35;
    sbox_4[51] = 8'd195;
    sbox_4[52] = 8'd24;
    sbox_4[53] = 8'd150;
    sbox_4[54] = 8'd5;
    sbox_4[55] = 8'd154;
    sbox_4[56] = 8'd7;
    sbox_4[57] = 8'd18;
    sbox_4[58] = 8'd128;
    sbox_4[59] = 8'd226;
    sbox_4[60] = 8'd235;
    sbox_4[61] = 8'd39;
    sbox_4[62] = 8'd178;
    sbox_4[63] = 8'd117;
    sbox_4[64] = 8'd9;
    sbox_4[65] = 8'd131;
    sbox_4[66] = 8'd44;
    sbox_4[67] = 8'd26;
    sbox_4[68] = 8'd27;
    sbox_4[69] = 8'd110;
    sbox_4[70] = 8'd90;
    sbox_4[71] = 8'd160;
    sbox_4[72] = 8'd82;
    sbox_4[73] = 8'd59;
    sbox_4[74] = 8'd214;
    sbox_4[75] = 8'd179;
    sbox_4[76] = 8'd41;
    sbox_4[77] = 8'd227;
    sbox_4[78] = 8'd47;
    sbox_4[79] = 8'd132;
    sbox_4[80] = 8'd83;
    sbox_4[81] = 8'd209;
    sbox_4[82] = 8'd0;
    sbox_4[83] = 8'd237;
    sbox_4[84] = 8'd32;
    sbox_4[85] = 8'd252;
    sbox_4[86] = 8'd177;
    sbox_4[87] = 8'd91;
    sbox_4[88] = 8'd106;
    sbox_4[89] = 8'd203;
    sbox_4[90] = 8'd190;
    sbox_4[91] = 8'd57;
    sbox_4[92] = 8'd74;
    sbox_4[93] = 8'd76;
    sbox_4[94] = 8'd88;
    sbox_4[95] = 8'd207;
    sbox_4[96] = 8'd208;
    sbox_4[97] = 8'd239;
    sbox_4[98] = 8'd170;
    sbox_4[99] = 8'd251;
    sbox_4[100] = 8'd67;
    sbox_4[101] = 8'd77;
    sbox_4[102] = 8'd51;
    sbox_4[103] = 8'd133;
    sbox_4[104] = 8'd69;
    sbox_4[105] = 8'd249;
    sbox_4[106] = 8'd2;
    sbox_4[107] = 8'd127;
    sbox_4[108] = 8'd80;
    sbox_4[109] = 8'd60;
    sbox_4[110] = 8'd159;
    sbox_4[111] = 8'd168;
    sbox_4[112] = 8'd81;
    sbox_4[113] = 8'd163;
    sbox_4[114] = 8'd64;
    sbox_4[115] = 8'd143;
    sbox_4[116] = 8'd146;
    sbox_4[117] = 8'd157;
    sbox_4[118] = 8'd56;
    sbox_4[119] = 8'd245;
    sbox_4[120] = 8'd188;
    sbox_4[121] = 8'd182;
    sbox_4[122] = 8'd218;
    sbox_4[123] = 8'd33;
    sbox_4[124] = 8'd16;
    sbox_4[125] = 8'd255;
    sbox_4[126] = 8'd243;
    sbox_4[127] = 8'd210;
    sbox_4[128] = 8'd205;
    sbox_4[129] = 8'd12;
    sbox_4[130] = 8'd19;
    sbox_4[131] = 8'd236;
    sbox_4[132] = 8'd95;
    sbox_4[133] = 8'd151;
    sbox_4[134] = 8'd68;
    sbox_4[135] = 8'd23;
    sbox_4[136] = 8'd196;
    sbox_4[137] = 8'd167;
    sbox_4[138] = 8'd126;
    sbox_4[139] = 8'd61;
    sbox_4[140] = 8'd100;
    sbox_4[141] = 8'd93;
    sbox_4[142] = 8'd25;
    sbox_4[143] = 8'd115;
    sbox_4[144] = 8'd96;
    sbox_4[145] = 8'd129;
    sbox_4[146] = 8'd79;
    sbox_4[147] = 8'd220;
    sbox_4[148] = 8'd34;
    sbox_4[149] = 8'd42;
    sbox_4[150] = 8'd144;
    sbox_4[151] = 8'd136;
    sbox_4[152] = 8'd70;
    sbox_4[153] = 8'd238;
    sbox_4[154] = 8'd184;
    sbox_4[155] = 8'd20;
    sbox_4[156] = 8'd222;
    sbox_4[157] = 8'd94;
    sbox_4[158] = 8'd11;
    sbox_4[159] = 8'd219;
    sbox_4[160] = 8'd224;
    sbox_4[161] = 8'd50;
    sbox_4[162] = 8'd58;
    sbox_4[163] = 8'd10;
    sbox_4[164] = 8'd73;
    sbox_4[165] = 8'd6;
    sbox_4[166] = 8'd36;
    sbox_4[167] = 8'd92;
    sbox_4[168] = 8'd194;
    sbox_4[169] = 8'd211;
    sbox_4[170] = 8'd172;
    sbox_4[171] = 8'd98;
    sbox_4[172] = 8'd145;
    sbox_4[173] = 8'd149;
    sbox_4[174] = 8'd228;
    sbox_4[175] = 8'd121;
    sbox_4[176] = 8'd231;
    sbox_4[177] = 8'd200;
    sbox_4[178] = 8'd55;
    sbox_4[179] = 8'd109;
    sbox_4[180] = 8'd141;
    sbox_4[181] = 8'd213;
    sbox_4[182] = 8'd78;
    sbox_4[183] = 8'd169;
    sbox_4[184] = 8'd108;
    sbox_4[185] = 8'd86;
    sbox_4[186] = 8'd244;
    sbox_4[187] = 8'd234;
    sbox_4[188] = 8'd101;
    sbox_4[189] = 8'd122;
    sbox_4[190] = 8'd174;
    sbox_4[191] = 8'd8;
    sbox_4[192] = 8'd186;
    sbox_4[193] = 8'd120;
    sbox_4[194] = 8'd37;
    sbox_4[195] = 8'd46;
    sbox_4[196] = 8'd28;
    sbox_4[197] = 8'd166;
    sbox_4[198] = 8'd180;
    sbox_4[199] = 8'd198;
    sbox_4[200] = 8'd232;
    sbox_4[201] = 8'd221;
    sbox_4[202] = 8'd116;
    sbox_4[203] = 8'd31;
    sbox_4[204] = 8'd75;
    sbox_4[205] = 8'd189;
    sbox_4[206] = 8'd139;
    sbox_4[207] = 8'd138;
    sbox_4[208] = 8'd112;
    sbox_4[209] = 8'd62;
    sbox_4[210] = 8'd181;
    sbox_4[211] = 8'd102;
    sbox_4[212] = 8'd72;
    sbox_4[213] = 8'd3;
    sbox_4[214] = 8'd246;
    sbox_4[215] = 8'd14;
    sbox_4[216] = 8'd97;
    sbox_4[217] = 8'd53;
    sbox_4[218] = 8'd87;
    sbox_4[219] = 8'd185;
    sbox_4[220] = 8'd134;
    sbox_4[221] = 8'd193;
    sbox_4[222] = 8'd29;
    sbox_4[223] = 8'd158;
    sbox_4[224] = 8'd225;
    sbox_4[225] = 8'd248;
    sbox_4[226] = 8'd152;
    sbox_4[227] = 8'd17;
    sbox_4[228] = 8'd105;
    sbox_4[229] = 8'd217;
    sbox_4[230] = 8'd142;
    sbox_4[231] = 8'd148;
    sbox_4[232] = 8'd155;
    sbox_4[233] = 8'd30;
    sbox_4[234] = 8'd135;
    sbox_4[235] = 8'd233;
    sbox_4[236] = 8'd206;
    sbox_4[237] = 8'd85;
    sbox_4[238] = 8'd40;
    sbox_4[239] = 8'd223;
    sbox_4[240] = 8'd140;
    sbox_4[241] = 8'd161;
    sbox_4[242] = 8'd137;
    sbox_4[243] = 8'd13;
    sbox_4[244] = 8'd191;
    sbox_4[245] = 8'd230;
    sbox_4[246] = 8'd66;
    sbox_4[247] = 8'd104;
    sbox_4[248] = 8'd65;
    sbox_4[249] = 8'd153;
    sbox_4[250] = 8'd45;
    sbox_4[251] = 8'd15;
    sbox_4[252] = 8'd176;
    sbox_4[253] = 8'd84;
    sbox_4[254] = 8'd187;
    sbox_4[255] = 8'd22;
    sbox_5[0] = 8'd99;
    sbox_5[1] = 8'd124;
    sbox_5[2] = 8'd119;
    sbox_5[3] = 8'd123;
    sbox_5[4] = 8'd242;
    sbox_5[5] = 8'd107;
    sbox_5[6] = 8'd111;
    sbox_5[7] = 8'd197;
    sbox_5[8] = 8'd48;
    sbox_5[9] = 8'd1;
    sbox_5[10] = 8'd103;
    sbox_5[11] = 8'd43;
    sbox_5[12] = 8'd254;
    sbox_5[13] = 8'd215;
    sbox_5[14] = 8'd171;
    sbox_5[15] = 8'd118;
    sbox_5[16] = 8'd202;
    sbox_5[17] = 8'd130;
    sbox_5[18] = 8'd201;
    sbox_5[19] = 8'd125;
    sbox_5[20] = 8'd250;
    sbox_5[21] = 8'd89;
    sbox_5[22] = 8'd71;
    sbox_5[23] = 8'd240;
    sbox_5[24] = 8'd173;
    sbox_5[25] = 8'd212;
    sbox_5[26] = 8'd162;
    sbox_5[27] = 8'd175;
    sbox_5[28] = 8'd156;
    sbox_5[29] = 8'd164;
    sbox_5[30] = 8'd114;
    sbox_5[31] = 8'd192;
    sbox_5[32] = 8'd183;
    sbox_5[33] = 8'd253;
    sbox_5[34] = 8'd147;
    sbox_5[35] = 8'd38;
    sbox_5[36] = 8'd54;
    sbox_5[37] = 8'd63;
    sbox_5[38] = 8'd247;
    sbox_5[39] = 8'd204;
    sbox_5[40] = 8'd52;
    sbox_5[41] = 8'd165;
    sbox_5[42] = 8'd229;
    sbox_5[43] = 8'd241;
    sbox_5[44] = 8'd113;
    sbox_5[45] = 8'd216;
    sbox_5[46] = 8'd49;
    sbox_5[47] = 8'd21;
    sbox_5[48] = 8'd4;
    sbox_5[49] = 8'd199;
    sbox_5[50] = 8'd35;
    sbox_5[51] = 8'd195;
    sbox_5[52] = 8'd24;
    sbox_5[53] = 8'd150;
    sbox_5[54] = 8'd5;
    sbox_5[55] = 8'd154;
    sbox_5[56] = 8'd7;
    sbox_5[57] = 8'd18;
    sbox_5[58] = 8'd128;
    sbox_5[59] = 8'd226;
    sbox_5[60] = 8'd235;
    sbox_5[61] = 8'd39;
    sbox_5[62] = 8'd178;
    sbox_5[63] = 8'd117;
    sbox_5[64] = 8'd9;
    sbox_5[65] = 8'd131;
    sbox_5[66] = 8'd44;
    sbox_5[67] = 8'd26;
    sbox_5[68] = 8'd27;
    sbox_5[69] = 8'd110;
    sbox_5[70] = 8'd90;
    sbox_5[71] = 8'd160;
    sbox_5[72] = 8'd82;
    sbox_5[73] = 8'd59;
    sbox_5[74] = 8'd214;
    sbox_5[75] = 8'd179;
    sbox_5[76] = 8'd41;
    sbox_5[77] = 8'd227;
    sbox_5[78] = 8'd47;
    sbox_5[79] = 8'd132;
    sbox_5[80] = 8'd83;
    sbox_5[81] = 8'd209;
    sbox_5[82] = 8'd0;
    sbox_5[83] = 8'd237;
    sbox_5[84] = 8'd32;
    sbox_5[85] = 8'd252;
    sbox_5[86] = 8'd177;
    sbox_5[87] = 8'd91;
    sbox_5[88] = 8'd106;
    sbox_5[89] = 8'd203;
    sbox_5[90] = 8'd190;
    sbox_5[91] = 8'd57;
    sbox_5[92] = 8'd74;
    sbox_5[93] = 8'd76;
    sbox_5[94] = 8'd88;
    sbox_5[95] = 8'd207;
    sbox_5[96] = 8'd208;
    sbox_5[97] = 8'd239;
    sbox_5[98] = 8'd170;
    sbox_5[99] = 8'd251;
    sbox_5[100] = 8'd67;
    sbox_5[101] = 8'd77;
    sbox_5[102] = 8'd51;
    sbox_5[103] = 8'd133;
    sbox_5[104] = 8'd69;
    sbox_5[105] = 8'd249;
    sbox_5[106] = 8'd2;
    sbox_5[107] = 8'd127;
    sbox_5[108] = 8'd80;
    sbox_5[109] = 8'd60;
    sbox_5[110] = 8'd159;
    sbox_5[111] = 8'd168;
    sbox_5[112] = 8'd81;
    sbox_5[113] = 8'd163;
    sbox_5[114] = 8'd64;
    sbox_5[115] = 8'd143;
    sbox_5[116] = 8'd146;
    sbox_5[117] = 8'd157;
    sbox_5[118] = 8'd56;
    sbox_5[119] = 8'd245;
    sbox_5[120] = 8'd188;
    sbox_5[121] = 8'd182;
    sbox_5[122] = 8'd218;
    sbox_5[123] = 8'd33;
    sbox_5[124] = 8'd16;
    sbox_5[125] = 8'd255;
    sbox_5[126] = 8'd243;
    sbox_5[127] = 8'd210;
    sbox_5[128] = 8'd205;
    sbox_5[129] = 8'd12;
    sbox_5[130] = 8'd19;
    sbox_5[131] = 8'd236;
    sbox_5[132] = 8'd95;
    sbox_5[133] = 8'd151;
    sbox_5[134] = 8'd68;
    sbox_5[135] = 8'd23;
    sbox_5[136] = 8'd196;
    sbox_5[137] = 8'd167;
    sbox_5[138] = 8'd126;
    sbox_5[139] = 8'd61;
    sbox_5[140] = 8'd100;
    sbox_5[141] = 8'd93;
    sbox_5[142] = 8'd25;
    sbox_5[143] = 8'd115;
    sbox_5[144] = 8'd96;
    sbox_5[145] = 8'd129;
    sbox_5[146] = 8'd79;
    sbox_5[147] = 8'd220;
    sbox_5[148] = 8'd34;
    sbox_5[149] = 8'd42;
    sbox_5[150] = 8'd144;
    sbox_5[151] = 8'd136;
    sbox_5[152] = 8'd70;
    sbox_5[153] = 8'd238;
    sbox_5[154] = 8'd184;
    sbox_5[155] = 8'd20;
    sbox_5[156] = 8'd222;
    sbox_5[157] = 8'd94;
    sbox_5[158] = 8'd11;
    sbox_5[159] = 8'd219;
    sbox_5[160] = 8'd224;
    sbox_5[161] = 8'd50;
    sbox_5[162] = 8'd58;
    sbox_5[163] = 8'd10;
    sbox_5[164] = 8'd73;
    sbox_5[165] = 8'd6;
    sbox_5[166] = 8'd36;
    sbox_5[167] = 8'd92;
    sbox_5[168] = 8'd194;
    sbox_5[169] = 8'd211;
    sbox_5[170] = 8'd172;
    sbox_5[171] = 8'd98;
    sbox_5[172] = 8'd145;
    sbox_5[173] = 8'd149;
    sbox_5[174] = 8'd228;
    sbox_5[175] = 8'd121;
    sbox_5[176] = 8'd231;
    sbox_5[177] = 8'd200;
    sbox_5[178] = 8'd55;
    sbox_5[179] = 8'd109;
    sbox_5[180] = 8'd141;
    sbox_5[181] = 8'd213;
    sbox_5[182] = 8'd78;
    sbox_5[183] = 8'd169;
    sbox_5[184] = 8'd108;
    sbox_5[185] = 8'd86;
    sbox_5[186] = 8'd244;
    sbox_5[187] = 8'd234;
    sbox_5[188] = 8'd101;
    sbox_5[189] = 8'd122;
    sbox_5[190] = 8'd174;
    sbox_5[191] = 8'd8;
    sbox_5[192] = 8'd186;
    sbox_5[193] = 8'd120;
    sbox_5[194] = 8'd37;
    sbox_5[195] = 8'd46;
    sbox_5[196] = 8'd28;
    sbox_5[197] = 8'd166;
    sbox_5[198] = 8'd180;
    sbox_5[199] = 8'd198;
    sbox_5[200] = 8'd232;
    sbox_5[201] = 8'd221;
    sbox_5[202] = 8'd116;
    sbox_5[203] = 8'd31;
    sbox_5[204] = 8'd75;
    sbox_5[205] = 8'd189;
    sbox_5[206] = 8'd139;
    sbox_5[207] = 8'd138;
    sbox_5[208] = 8'd112;
    sbox_5[209] = 8'd62;
    sbox_5[210] = 8'd181;
    sbox_5[211] = 8'd102;
    sbox_5[212] = 8'd72;
    sbox_5[213] = 8'd3;
    sbox_5[214] = 8'd246;
    sbox_5[215] = 8'd14;
    sbox_5[216] = 8'd97;
    sbox_5[217] = 8'd53;
    sbox_5[218] = 8'd87;
    sbox_5[219] = 8'd185;
    sbox_5[220] = 8'd134;
    sbox_5[221] = 8'd193;
    sbox_5[222] = 8'd29;
    sbox_5[223] = 8'd158;
    sbox_5[224] = 8'd225;
    sbox_5[225] = 8'd248;
    sbox_5[226] = 8'd152;
    sbox_5[227] = 8'd17;
    sbox_5[228] = 8'd105;
    sbox_5[229] = 8'd217;
    sbox_5[230] = 8'd142;
    sbox_5[231] = 8'd148;
    sbox_5[232] = 8'd155;
    sbox_5[233] = 8'd30;
    sbox_5[234] = 8'd135;
    sbox_5[235] = 8'd233;
    sbox_5[236] = 8'd206;
    sbox_5[237] = 8'd85;
    sbox_5[238] = 8'd40;
    sbox_5[239] = 8'd223;
    sbox_5[240] = 8'd140;
    sbox_5[241] = 8'd161;
    sbox_5[242] = 8'd137;
    sbox_5[243] = 8'd13;
    sbox_5[244] = 8'd191;
    sbox_5[245] = 8'd230;
    sbox_5[246] = 8'd66;
    sbox_5[247] = 8'd104;
    sbox_5[248] = 8'd65;
    sbox_5[249] = 8'd153;
    sbox_5[250] = 8'd45;
    sbox_5[251] = 8'd15;
    sbox_5[252] = 8'd176;
    sbox_5[253] = 8'd84;
    sbox_5[254] = 8'd187;
    sbox_5[255] = 8'd22;
    sbox_6[0] = 8'd99;
    sbox_6[1] = 8'd124;
    sbox_6[2] = 8'd119;
    sbox_6[3] = 8'd123;
    sbox_6[4] = 8'd242;
    sbox_6[5] = 8'd107;
    sbox_6[6] = 8'd111;
    sbox_6[7] = 8'd197;
    sbox_6[8] = 8'd48;
    sbox_6[9] = 8'd1;
    sbox_6[10] = 8'd103;
    sbox_6[11] = 8'd43;
    sbox_6[12] = 8'd254;
    sbox_6[13] = 8'd215;
    sbox_6[14] = 8'd171;
    sbox_6[15] = 8'd118;
    sbox_6[16] = 8'd202;
    sbox_6[17] = 8'd130;
    sbox_6[18] = 8'd201;
    sbox_6[19] = 8'd125;
    sbox_6[20] = 8'd250;
    sbox_6[21] = 8'd89;
    sbox_6[22] = 8'd71;
    sbox_6[23] = 8'd240;
    sbox_6[24] = 8'd173;
    sbox_6[25] = 8'd212;
    sbox_6[26] = 8'd162;
    sbox_6[27] = 8'd175;
    sbox_6[28] = 8'd156;
    sbox_6[29] = 8'd164;
    sbox_6[30] = 8'd114;
    sbox_6[31] = 8'd192;
    sbox_6[32] = 8'd183;
    sbox_6[33] = 8'd253;
    sbox_6[34] = 8'd147;
    sbox_6[35] = 8'd38;
    sbox_6[36] = 8'd54;
    sbox_6[37] = 8'd63;
    sbox_6[38] = 8'd247;
    sbox_6[39] = 8'd204;
    sbox_6[40] = 8'd52;
    sbox_6[41] = 8'd165;
    sbox_6[42] = 8'd229;
    sbox_6[43] = 8'd241;
    sbox_6[44] = 8'd113;
    sbox_6[45] = 8'd216;
    sbox_6[46] = 8'd49;
    sbox_6[47] = 8'd21;
    sbox_6[48] = 8'd4;
    sbox_6[49] = 8'd199;
    sbox_6[50] = 8'd35;
    sbox_6[51] = 8'd195;
    sbox_6[52] = 8'd24;
    sbox_6[53] = 8'd150;
    sbox_6[54] = 8'd5;
    sbox_6[55] = 8'd154;
    sbox_6[56] = 8'd7;
    sbox_6[57] = 8'd18;
    sbox_6[58] = 8'd128;
    sbox_6[59] = 8'd226;
    sbox_6[60] = 8'd235;
    sbox_6[61] = 8'd39;
    sbox_6[62] = 8'd178;
    sbox_6[63] = 8'd117;
    sbox_6[64] = 8'd9;
    sbox_6[65] = 8'd131;
    sbox_6[66] = 8'd44;
    sbox_6[67] = 8'd26;
    sbox_6[68] = 8'd27;
    sbox_6[69] = 8'd110;
    sbox_6[70] = 8'd90;
    sbox_6[71] = 8'd160;
    sbox_6[72] = 8'd82;
    sbox_6[73] = 8'd59;
    sbox_6[74] = 8'd214;
    sbox_6[75] = 8'd179;
    sbox_6[76] = 8'd41;
    sbox_6[77] = 8'd227;
    sbox_6[78] = 8'd47;
    sbox_6[79] = 8'd132;
    sbox_6[80] = 8'd83;
    sbox_6[81] = 8'd209;
    sbox_6[82] = 8'd0;
    sbox_6[83] = 8'd237;
    sbox_6[84] = 8'd32;
    sbox_6[85] = 8'd252;
    sbox_6[86] = 8'd177;
    sbox_6[87] = 8'd91;
    sbox_6[88] = 8'd106;
    sbox_6[89] = 8'd203;
    sbox_6[90] = 8'd190;
    sbox_6[91] = 8'd57;
    sbox_6[92] = 8'd74;
    sbox_6[93] = 8'd76;
    sbox_6[94] = 8'd88;
    sbox_6[95] = 8'd207;
    sbox_6[96] = 8'd208;
    sbox_6[97] = 8'd239;
    sbox_6[98] = 8'd170;
    sbox_6[99] = 8'd251;
    sbox_6[100] = 8'd67;
    sbox_6[101] = 8'd77;
    sbox_6[102] = 8'd51;
    sbox_6[103] = 8'd133;
    sbox_6[104] = 8'd69;
    sbox_6[105] = 8'd249;
    sbox_6[106] = 8'd2;
    sbox_6[107] = 8'd127;
    sbox_6[108] = 8'd80;
    sbox_6[109] = 8'd60;
    sbox_6[110] = 8'd159;
    sbox_6[111] = 8'd168;
    sbox_6[112] = 8'd81;
    sbox_6[113] = 8'd163;
    sbox_6[114] = 8'd64;
    sbox_6[115] = 8'd143;
    sbox_6[116] = 8'd146;
    sbox_6[117] = 8'd157;
    sbox_6[118] = 8'd56;
    sbox_6[119] = 8'd245;
    sbox_6[120] = 8'd188;
    sbox_6[121] = 8'd182;
    sbox_6[122] = 8'd218;
    sbox_6[123] = 8'd33;
    sbox_6[124] = 8'd16;
    sbox_6[125] = 8'd255;
    sbox_6[126] = 8'd243;
    sbox_6[127] = 8'd210;
    sbox_6[128] = 8'd205;
    sbox_6[129] = 8'd12;
    sbox_6[130] = 8'd19;
    sbox_6[131] = 8'd236;
    sbox_6[132] = 8'd95;
    sbox_6[133] = 8'd151;
    sbox_6[134] = 8'd68;
    sbox_6[135] = 8'd23;
    sbox_6[136] = 8'd196;
    sbox_6[137] = 8'd167;
    sbox_6[138] = 8'd126;
    sbox_6[139] = 8'd61;
    sbox_6[140] = 8'd100;
    sbox_6[141] = 8'd93;
    sbox_6[142] = 8'd25;
    sbox_6[143] = 8'd115;
    sbox_6[144] = 8'd96;
    sbox_6[145] = 8'd129;
    sbox_6[146] = 8'd79;
    sbox_6[147] = 8'd220;
    sbox_6[148] = 8'd34;
    sbox_6[149] = 8'd42;
    sbox_6[150] = 8'd144;
    sbox_6[151] = 8'd136;
    sbox_6[152] = 8'd70;
    sbox_6[153] = 8'd238;
    sbox_6[154] = 8'd184;
    sbox_6[155] = 8'd20;
    sbox_6[156] = 8'd222;
    sbox_6[157] = 8'd94;
    sbox_6[158] = 8'd11;
    sbox_6[159] = 8'd219;
    sbox_6[160] = 8'd224;
    sbox_6[161] = 8'd50;
    sbox_6[162] = 8'd58;
    sbox_6[163] = 8'd10;
    sbox_6[164] = 8'd73;
    sbox_6[165] = 8'd6;
    sbox_6[166] = 8'd36;
    sbox_6[167] = 8'd92;
    sbox_6[168] = 8'd194;
    sbox_6[169] = 8'd211;
    sbox_6[170] = 8'd172;
    sbox_6[171] = 8'd98;
    sbox_6[172] = 8'd145;
    sbox_6[173] = 8'd149;
    sbox_6[174] = 8'd228;
    sbox_6[175] = 8'd121;
    sbox_6[176] = 8'd231;
    sbox_6[177] = 8'd200;
    sbox_6[178] = 8'd55;
    sbox_6[179] = 8'd109;
    sbox_6[180] = 8'd141;
    sbox_6[181] = 8'd213;
    sbox_6[182] = 8'd78;
    sbox_6[183] = 8'd169;
    sbox_6[184] = 8'd108;
    sbox_6[185] = 8'd86;
    sbox_6[186] = 8'd244;
    sbox_6[187] = 8'd234;
    sbox_6[188] = 8'd101;
    sbox_6[189] = 8'd122;
    sbox_6[190] = 8'd174;
    sbox_6[191] = 8'd8;
    sbox_6[192] = 8'd186;
    sbox_6[193] = 8'd120;
    sbox_6[194] = 8'd37;
    sbox_6[195] = 8'd46;
    sbox_6[196] = 8'd28;
    sbox_6[197] = 8'd166;
    sbox_6[198] = 8'd180;
    sbox_6[199] = 8'd198;
    sbox_6[200] = 8'd232;
    sbox_6[201] = 8'd221;
    sbox_6[202] = 8'd116;
    sbox_6[203] = 8'd31;
    sbox_6[204] = 8'd75;
    sbox_6[205] = 8'd189;
    sbox_6[206] = 8'd139;
    sbox_6[207] = 8'd138;
    sbox_6[208] = 8'd112;
    sbox_6[209] = 8'd62;
    sbox_6[210] = 8'd181;
    sbox_6[211] = 8'd102;
    sbox_6[212] = 8'd72;
    sbox_6[213] = 8'd3;
    sbox_6[214] = 8'd246;
    sbox_6[215] = 8'd14;
    sbox_6[216] = 8'd97;
    sbox_6[217] = 8'd53;
    sbox_6[218] = 8'd87;
    sbox_6[219] = 8'd185;
    sbox_6[220] = 8'd134;
    sbox_6[221] = 8'd193;
    sbox_6[222] = 8'd29;
    sbox_6[223] = 8'd158;
    sbox_6[224] = 8'd225;
    sbox_6[225] = 8'd248;
    sbox_6[226] = 8'd152;
    sbox_6[227] = 8'd17;
    sbox_6[228] = 8'd105;
    sbox_6[229] = 8'd217;
    sbox_6[230] = 8'd142;
    sbox_6[231] = 8'd148;
    sbox_6[232] = 8'd155;
    sbox_6[233] = 8'd30;
    sbox_6[234] = 8'd135;
    sbox_6[235] = 8'd233;
    sbox_6[236] = 8'd206;
    sbox_6[237] = 8'd85;
    sbox_6[238] = 8'd40;
    sbox_6[239] = 8'd223;
    sbox_6[240] = 8'd140;
    sbox_6[241] = 8'd161;
    sbox_6[242] = 8'd137;
    sbox_6[243] = 8'd13;
    sbox_6[244] = 8'd191;
    sbox_6[245] = 8'd230;
    sbox_6[246] = 8'd66;
    sbox_6[247] = 8'd104;
    sbox_6[248] = 8'd65;
    sbox_6[249] = 8'd153;
    sbox_6[250] = 8'd45;
    sbox_6[251] = 8'd15;
    sbox_6[252] = 8'd176;
    sbox_6[253] = 8'd84;
    sbox_6[254] = 8'd187;
    sbox_6[255] = 8'd22;
    sbox_7[0] = 8'd99;
    sbox_7[1] = 8'd124;
    sbox_7[2] = 8'd119;
    sbox_7[3] = 8'd123;
    sbox_7[4] = 8'd242;
    sbox_7[5] = 8'd107;
    sbox_7[6] = 8'd111;
    sbox_7[7] = 8'd197;
    sbox_7[8] = 8'd48;
    sbox_7[9] = 8'd1;
    sbox_7[10] = 8'd103;
    sbox_7[11] = 8'd43;
    sbox_7[12] = 8'd254;
    sbox_7[13] = 8'd215;
    sbox_7[14] = 8'd171;
    sbox_7[15] = 8'd118;
    sbox_7[16] = 8'd202;
    sbox_7[17] = 8'd130;
    sbox_7[18] = 8'd201;
    sbox_7[19] = 8'd125;
    sbox_7[20] = 8'd250;
    sbox_7[21] = 8'd89;
    sbox_7[22] = 8'd71;
    sbox_7[23] = 8'd240;
    sbox_7[24] = 8'd173;
    sbox_7[25] = 8'd212;
    sbox_7[26] = 8'd162;
    sbox_7[27] = 8'd175;
    sbox_7[28] = 8'd156;
    sbox_7[29] = 8'd164;
    sbox_7[30] = 8'd114;
    sbox_7[31] = 8'd192;
    sbox_7[32] = 8'd183;
    sbox_7[33] = 8'd253;
    sbox_7[34] = 8'd147;
    sbox_7[35] = 8'd38;
    sbox_7[36] = 8'd54;
    sbox_7[37] = 8'd63;
    sbox_7[38] = 8'd247;
    sbox_7[39] = 8'd204;
    sbox_7[40] = 8'd52;
    sbox_7[41] = 8'd165;
    sbox_7[42] = 8'd229;
    sbox_7[43] = 8'd241;
    sbox_7[44] = 8'd113;
    sbox_7[45] = 8'd216;
    sbox_7[46] = 8'd49;
    sbox_7[47] = 8'd21;
    sbox_7[48] = 8'd4;
    sbox_7[49] = 8'd199;
    sbox_7[50] = 8'd35;
    sbox_7[51] = 8'd195;
    sbox_7[52] = 8'd24;
    sbox_7[53] = 8'd150;
    sbox_7[54] = 8'd5;
    sbox_7[55] = 8'd154;
    sbox_7[56] = 8'd7;
    sbox_7[57] = 8'd18;
    sbox_7[58] = 8'd128;
    sbox_7[59] = 8'd226;
    sbox_7[60] = 8'd235;
    sbox_7[61] = 8'd39;
    sbox_7[62] = 8'd178;
    sbox_7[63] = 8'd117;
    sbox_7[64] = 8'd9;
    sbox_7[65] = 8'd131;
    sbox_7[66] = 8'd44;
    sbox_7[67] = 8'd26;
    sbox_7[68] = 8'd27;
    sbox_7[69] = 8'd110;
    sbox_7[70] = 8'd90;
    sbox_7[71] = 8'd160;
    sbox_7[72] = 8'd82;
    sbox_7[73] = 8'd59;
    sbox_7[74] = 8'd214;
    sbox_7[75] = 8'd179;
    sbox_7[76] = 8'd41;
    sbox_7[77] = 8'd227;
    sbox_7[78] = 8'd47;
    sbox_7[79] = 8'd132;
    sbox_7[80] = 8'd83;
    sbox_7[81] = 8'd209;
    sbox_7[82] = 8'd0;
    sbox_7[83] = 8'd237;
    sbox_7[84] = 8'd32;
    sbox_7[85] = 8'd252;
    sbox_7[86] = 8'd177;
    sbox_7[87] = 8'd91;
    sbox_7[88] = 8'd106;
    sbox_7[89] = 8'd203;
    sbox_7[90] = 8'd190;
    sbox_7[91] = 8'd57;
    sbox_7[92] = 8'd74;
    sbox_7[93] = 8'd76;
    sbox_7[94] = 8'd88;
    sbox_7[95] = 8'd207;
    sbox_7[96] = 8'd208;
    sbox_7[97] = 8'd239;
    sbox_7[98] = 8'd170;
    sbox_7[99] = 8'd251;
    sbox_7[100] = 8'd67;
    sbox_7[101] = 8'd77;
    sbox_7[102] = 8'd51;
    sbox_7[103] = 8'd133;
    sbox_7[104] = 8'd69;
    sbox_7[105] = 8'd249;
    sbox_7[106] = 8'd2;
    sbox_7[107] = 8'd127;
    sbox_7[108] = 8'd80;
    sbox_7[109] = 8'd60;
    sbox_7[110] = 8'd159;
    sbox_7[111] = 8'd168;
    sbox_7[112] = 8'd81;
    sbox_7[113] = 8'd163;
    sbox_7[114] = 8'd64;
    sbox_7[115] = 8'd143;
    sbox_7[116] = 8'd146;
    sbox_7[117] = 8'd157;
    sbox_7[118] = 8'd56;
    sbox_7[119] = 8'd245;
    sbox_7[120] = 8'd188;
    sbox_7[121] = 8'd182;
    sbox_7[122] = 8'd218;
    sbox_7[123] = 8'd33;
    sbox_7[124] = 8'd16;
    sbox_7[125] = 8'd255;
    sbox_7[126] = 8'd243;
    sbox_7[127] = 8'd210;
    sbox_7[128] = 8'd205;
    sbox_7[129] = 8'd12;
    sbox_7[130] = 8'd19;
    sbox_7[131] = 8'd236;
    sbox_7[132] = 8'd95;
    sbox_7[133] = 8'd151;
    sbox_7[134] = 8'd68;
    sbox_7[135] = 8'd23;
    sbox_7[136] = 8'd196;
    sbox_7[137] = 8'd167;
    sbox_7[138] = 8'd126;
    sbox_7[139] = 8'd61;
    sbox_7[140] = 8'd100;
    sbox_7[141] = 8'd93;
    sbox_7[142] = 8'd25;
    sbox_7[143] = 8'd115;
    sbox_7[144] = 8'd96;
    sbox_7[145] = 8'd129;
    sbox_7[146] = 8'd79;
    sbox_7[147] = 8'd220;
    sbox_7[148] = 8'd34;
    sbox_7[149] = 8'd42;
    sbox_7[150] = 8'd144;
    sbox_7[151] = 8'd136;
    sbox_7[152] = 8'd70;
    sbox_7[153] = 8'd238;
    sbox_7[154] = 8'd184;
    sbox_7[155] = 8'd20;
    sbox_7[156] = 8'd222;
    sbox_7[157] = 8'd94;
    sbox_7[158] = 8'd11;
    sbox_7[159] = 8'd219;
    sbox_7[160] = 8'd224;
    sbox_7[161] = 8'd50;
    sbox_7[162] = 8'd58;
    sbox_7[163] = 8'd10;
    sbox_7[164] = 8'd73;
    sbox_7[165] = 8'd6;
    sbox_7[166] = 8'd36;
    sbox_7[167] = 8'd92;
    sbox_7[168] = 8'd194;
    sbox_7[169] = 8'd211;
    sbox_7[170] = 8'd172;
    sbox_7[171] = 8'd98;
    sbox_7[172] = 8'd145;
    sbox_7[173] = 8'd149;
    sbox_7[174] = 8'd228;
    sbox_7[175] = 8'd121;
    sbox_7[176] = 8'd231;
    sbox_7[177] = 8'd200;
    sbox_7[178] = 8'd55;
    sbox_7[179] = 8'd109;
    sbox_7[180] = 8'd141;
    sbox_7[181] = 8'd213;
    sbox_7[182] = 8'd78;
    sbox_7[183] = 8'd169;
    sbox_7[184] = 8'd108;
    sbox_7[185] = 8'd86;
    sbox_7[186] = 8'd244;
    sbox_7[187] = 8'd234;
    sbox_7[188] = 8'd101;
    sbox_7[189] = 8'd122;
    sbox_7[190] = 8'd174;
    sbox_7[191] = 8'd8;
    sbox_7[192] = 8'd186;
    sbox_7[193] = 8'd120;
    sbox_7[194] = 8'd37;
    sbox_7[195] = 8'd46;
    sbox_7[196] = 8'd28;
    sbox_7[197] = 8'd166;
    sbox_7[198] = 8'd180;
    sbox_7[199] = 8'd198;
    sbox_7[200] = 8'd232;
    sbox_7[201] = 8'd221;
    sbox_7[202] = 8'd116;
    sbox_7[203] = 8'd31;
    sbox_7[204] = 8'd75;
    sbox_7[205] = 8'd189;
    sbox_7[206] = 8'd139;
    sbox_7[207] = 8'd138;
    sbox_7[208] = 8'd112;
    sbox_7[209] = 8'd62;
    sbox_7[210] = 8'd181;
    sbox_7[211] = 8'd102;
    sbox_7[212] = 8'd72;
    sbox_7[213] = 8'd3;
    sbox_7[214] = 8'd246;
    sbox_7[215] = 8'd14;
    sbox_7[216] = 8'd97;
    sbox_7[217] = 8'd53;
    sbox_7[218] = 8'd87;
    sbox_7[219] = 8'd185;
    sbox_7[220] = 8'd134;
    sbox_7[221] = 8'd193;
    sbox_7[222] = 8'd29;
    sbox_7[223] = 8'd158;
    sbox_7[224] = 8'd225;
    sbox_7[225] = 8'd248;
    sbox_7[226] = 8'd152;
    sbox_7[227] = 8'd17;
    sbox_7[228] = 8'd105;
    sbox_7[229] = 8'd217;
    sbox_7[230] = 8'd142;
    sbox_7[231] = 8'd148;
    sbox_7[232] = 8'd155;
    sbox_7[233] = 8'd30;
    sbox_7[234] = 8'd135;
    sbox_7[235] = 8'd233;
    sbox_7[236] = 8'd206;
    sbox_7[237] = 8'd85;
    sbox_7[238] = 8'd40;
    sbox_7[239] = 8'd223;
    sbox_7[240] = 8'd140;
    sbox_7[241] = 8'd161;
    sbox_7[242] = 8'd137;
    sbox_7[243] = 8'd13;
    sbox_7[244] = 8'd191;
    sbox_7[245] = 8'd230;
    sbox_7[246] = 8'd66;
    sbox_7[247] = 8'd104;
    sbox_7[248] = 8'd65;
    sbox_7[249] = 8'd153;
    sbox_7[250] = 8'd45;
    sbox_7[251] = 8'd15;
    sbox_7[252] = 8'd176;
    sbox_7[253] = 8'd84;
    sbox_7[254] = 8'd187;
    sbox_7[255] = 8'd22;
    sbox_8[0] = 8'd99;
    sbox_8[1] = 8'd124;
    sbox_8[2] = 8'd119;
    sbox_8[3] = 8'd123;
    sbox_8[4] = 8'd242;
    sbox_8[5] = 8'd107;
    sbox_8[6] = 8'd111;
    sbox_8[7] = 8'd197;
    sbox_8[8] = 8'd48;
    sbox_8[9] = 8'd1;
    sbox_8[10] = 8'd103;
    sbox_8[11] = 8'd43;
    sbox_8[12] = 8'd254;
    sbox_8[13] = 8'd215;
    sbox_8[14] = 8'd171;
    sbox_8[15] = 8'd118;
    sbox_8[16] = 8'd202;
    sbox_8[17] = 8'd130;
    sbox_8[18] = 8'd201;
    sbox_8[19] = 8'd125;
    sbox_8[20] = 8'd250;
    sbox_8[21] = 8'd89;
    sbox_8[22] = 8'd71;
    sbox_8[23] = 8'd240;
    sbox_8[24] = 8'd173;
    sbox_8[25] = 8'd212;
    sbox_8[26] = 8'd162;
    sbox_8[27] = 8'd175;
    sbox_8[28] = 8'd156;
    sbox_8[29] = 8'd164;
    sbox_8[30] = 8'd114;
    sbox_8[31] = 8'd192;
    sbox_8[32] = 8'd183;
    sbox_8[33] = 8'd253;
    sbox_8[34] = 8'd147;
    sbox_8[35] = 8'd38;
    sbox_8[36] = 8'd54;
    sbox_8[37] = 8'd63;
    sbox_8[38] = 8'd247;
    sbox_8[39] = 8'd204;
    sbox_8[40] = 8'd52;
    sbox_8[41] = 8'd165;
    sbox_8[42] = 8'd229;
    sbox_8[43] = 8'd241;
    sbox_8[44] = 8'd113;
    sbox_8[45] = 8'd216;
    sbox_8[46] = 8'd49;
    sbox_8[47] = 8'd21;
    sbox_8[48] = 8'd4;
    sbox_8[49] = 8'd199;
    sbox_8[50] = 8'd35;
    sbox_8[51] = 8'd195;
    sbox_8[52] = 8'd24;
    sbox_8[53] = 8'd150;
    sbox_8[54] = 8'd5;
    sbox_8[55] = 8'd154;
    sbox_8[56] = 8'd7;
    sbox_8[57] = 8'd18;
    sbox_8[58] = 8'd128;
    sbox_8[59] = 8'd226;
    sbox_8[60] = 8'd235;
    sbox_8[61] = 8'd39;
    sbox_8[62] = 8'd178;
    sbox_8[63] = 8'd117;
    sbox_8[64] = 8'd9;
    sbox_8[65] = 8'd131;
    sbox_8[66] = 8'd44;
    sbox_8[67] = 8'd26;
    sbox_8[68] = 8'd27;
    sbox_8[69] = 8'd110;
    sbox_8[70] = 8'd90;
    sbox_8[71] = 8'd160;
    sbox_8[72] = 8'd82;
    sbox_8[73] = 8'd59;
    sbox_8[74] = 8'd214;
    sbox_8[75] = 8'd179;
    sbox_8[76] = 8'd41;
    sbox_8[77] = 8'd227;
    sbox_8[78] = 8'd47;
    sbox_8[79] = 8'd132;
    sbox_8[80] = 8'd83;
    sbox_8[81] = 8'd209;
    sbox_8[82] = 8'd0;
    sbox_8[83] = 8'd237;
    sbox_8[84] = 8'd32;
    sbox_8[85] = 8'd252;
    sbox_8[86] = 8'd177;
    sbox_8[87] = 8'd91;
    sbox_8[88] = 8'd106;
    sbox_8[89] = 8'd203;
    sbox_8[90] = 8'd190;
    sbox_8[91] = 8'd57;
    sbox_8[92] = 8'd74;
    sbox_8[93] = 8'd76;
    sbox_8[94] = 8'd88;
    sbox_8[95] = 8'd207;
    sbox_8[96] = 8'd208;
    sbox_8[97] = 8'd239;
    sbox_8[98] = 8'd170;
    sbox_8[99] = 8'd251;
    sbox_8[100] = 8'd67;
    sbox_8[101] = 8'd77;
    sbox_8[102] = 8'd51;
    sbox_8[103] = 8'd133;
    sbox_8[104] = 8'd69;
    sbox_8[105] = 8'd249;
    sbox_8[106] = 8'd2;
    sbox_8[107] = 8'd127;
    sbox_8[108] = 8'd80;
    sbox_8[109] = 8'd60;
    sbox_8[110] = 8'd159;
    sbox_8[111] = 8'd168;
    sbox_8[112] = 8'd81;
    sbox_8[113] = 8'd163;
    sbox_8[114] = 8'd64;
    sbox_8[115] = 8'd143;
    sbox_8[116] = 8'd146;
    sbox_8[117] = 8'd157;
    sbox_8[118] = 8'd56;
    sbox_8[119] = 8'd245;
    sbox_8[120] = 8'd188;
    sbox_8[121] = 8'd182;
    sbox_8[122] = 8'd218;
    sbox_8[123] = 8'd33;
    sbox_8[124] = 8'd16;
    sbox_8[125] = 8'd255;
    sbox_8[126] = 8'd243;
    sbox_8[127] = 8'd210;
    sbox_8[128] = 8'd205;
    sbox_8[129] = 8'd12;
    sbox_8[130] = 8'd19;
    sbox_8[131] = 8'd236;
    sbox_8[132] = 8'd95;
    sbox_8[133] = 8'd151;
    sbox_8[134] = 8'd68;
    sbox_8[135] = 8'd23;
    sbox_8[136] = 8'd196;
    sbox_8[137] = 8'd167;
    sbox_8[138] = 8'd126;
    sbox_8[139] = 8'd61;
    sbox_8[140] = 8'd100;
    sbox_8[141] = 8'd93;
    sbox_8[142] = 8'd25;
    sbox_8[143] = 8'd115;
    sbox_8[144] = 8'd96;
    sbox_8[145] = 8'd129;
    sbox_8[146] = 8'd79;
    sbox_8[147] = 8'd220;
    sbox_8[148] = 8'd34;
    sbox_8[149] = 8'd42;
    sbox_8[150] = 8'd144;
    sbox_8[151] = 8'd136;
    sbox_8[152] = 8'd70;
    sbox_8[153] = 8'd238;
    sbox_8[154] = 8'd184;
    sbox_8[155] = 8'd20;
    sbox_8[156] = 8'd222;
    sbox_8[157] = 8'd94;
    sbox_8[158] = 8'd11;
    sbox_8[159] = 8'd219;
    sbox_8[160] = 8'd224;
    sbox_8[161] = 8'd50;
    sbox_8[162] = 8'd58;
    sbox_8[163] = 8'd10;
    sbox_8[164] = 8'd73;
    sbox_8[165] = 8'd6;
    sbox_8[166] = 8'd36;
    sbox_8[167] = 8'd92;
    sbox_8[168] = 8'd194;
    sbox_8[169] = 8'd211;
    sbox_8[170] = 8'd172;
    sbox_8[171] = 8'd98;
    sbox_8[172] = 8'd145;
    sbox_8[173] = 8'd149;
    sbox_8[174] = 8'd228;
    sbox_8[175] = 8'd121;
    sbox_8[176] = 8'd231;
    sbox_8[177] = 8'd200;
    sbox_8[178] = 8'd55;
    sbox_8[179] = 8'd109;
    sbox_8[180] = 8'd141;
    sbox_8[181] = 8'd213;
    sbox_8[182] = 8'd78;
    sbox_8[183] = 8'd169;
    sbox_8[184] = 8'd108;
    sbox_8[185] = 8'd86;
    sbox_8[186] = 8'd244;
    sbox_8[187] = 8'd234;
    sbox_8[188] = 8'd101;
    sbox_8[189] = 8'd122;
    sbox_8[190] = 8'd174;
    sbox_8[191] = 8'd8;
    sbox_8[192] = 8'd186;
    sbox_8[193] = 8'd120;
    sbox_8[194] = 8'd37;
    sbox_8[195] = 8'd46;
    sbox_8[196] = 8'd28;
    sbox_8[197] = 8'd166;
    sbox_8[198] = 8'd180;
    sbox_8[199] = 8'd198;
    sbox_8[200] = 8'd232;
    sbox_8[201] = 8'd221;
    sbox_8[202] = 8'd116;
    sbox_8[203] = 8'd31;
    sbox_8[204] = 8'd75;
    sbox_8[205] = 8'd189;
    sbox_8[206] = 8'd139;
    sbox_8[207] = 8'd138;
    sbox_8[208] = 8'd112;
    sbox_8[209] = 8'd62;
    sbox_8[210] = 8'd181;
    sbox_8[211] = 8'd102;
    sbox_8[212] = 8'd72;
    sbox_8[213] = 8'd3;
    sbox_8[214] = 8'd246;
    sbox_8[215] = 8'd14;
    sbox_8[216] = 8'd97;
    sbox_8[217] = 8'd53;
    sbox_8[218] = 8'd87;
    sbox_8[219] = 8'd185;
    sbox_8[220] = 8'd134;
    sbox_8[221] = 8'd193;
    sbox_8[222] = 8'd29;
    sbox_8[223] = 8'd158;
    sbox_8[224] = 8'd225;
    sbox_8[225] = 8'd248;
    sbox_8[226] = 8'd152;
    sbox_8[227] = 8'd17;
    sbox_8[228] = 8'd105;
    sbox_8[229] = 8'd217;
    sbox_8[230] = 8'd142;
    sbox_8[231] = 8'd148;
    sbox_8[232] = 8'd155;
    sbox_8[233] = 8'd30;
    sbox_8[234] = 8'd135;
    sbox_8[235] = 8'd233;
    sbox_8[236] = 8'd206;
    sbox_8[237] = 8'd85;
    sbox_8[238] = 8'd40;
    sbox_8[239] = 8'd223;
    sbox_8[240] = 8'd140;
    sbox_8[241] = 8'd161;
    sbox_8[242] = 8'd137;
    sbox_8[243] = 8'd13;
    sbox_8[244] = 8'd191;
    sbox_8[245] = 8'd230;
    sbox_8[246] = 8'd66;
    sbox_8[247] = 8'd104;
    sbox_8[248] = 8'd65;
    sbox_8[249] = 8'd153;
    sbox_8[250] = 8'd45;
    sbox_8[251] = 8'd15;
    sbox_8[252] = 8'd176;
    sbox_8[253] = 8'd84;
    sbox_8[254] = 8'd187;
    sbox_8[255] = 8'd22;
    sbox_9[0] = 8'd99;
    sbox_9[1] = 8'd124;
    sbox_9[2] = 8'd119;
    sbox_9[3] = 8'd123;
    sbox_9[4] = 8'd242;
    sbox_9[5] = 8'd107;
    sbox_9[6] = 8'd111;
    sbox_9[7] = 8'd197;
    sbox_9[8] = 8'd48;
    sbox_9[9] = 8'd1;
    sbox_9[10] = 8'd103;
    sbox_9[11] = 8'd43;
    sbox_9[12] = 8'd254;
    sbox_9[13] = 8'd215;
    sbox_9[14] = 8'd171;
    sbox_9[15] = 8'd118;
    sbox_9[16] = 8'd202;
    sbox_9[17] = 8'd130;
    sbox_9[18] = 8'd201;
    sbox_9[19] = 8'd125;
    sbox_9[20] = 8'd250;
    sbox_9[21] = 8'd89;
    sbox_9[22] = 8'd71;
    sbox_9[23] = 8'd240;
    sbox_9[24] = 8'd173;
    sbox_9[25] = 8'd212;
    sbox_9[26] = 8'd162;
    sbox_9[27] = 8'd175;
    sbox_9[28] = 8'd156;
    sbox_9[29] = 8'd164;
    sbox_9[30] = 8'd114;
    sbox_9[31] = 8'd192;
    sbox_9[32] = 8'd183;
    sbox_9[33] = 8'd253;
    sbox_9[34] = 8'd147;
    sbox_9[35] = 8'd38;
    sbox_9[36] = 8'd54;
    sbox_9[37] = 8'd63;
    sbox_9[38] = 8'd247;
    sbox_9[39] = 8'd204;
    sbox_9[40] = 8'd52;
    sbox_9[41] = 8'd165;
    sbox_9[42] = 8'd229;
    sbox_9[43] = 8'd241;
    sbox_9[44] = 8'd113;
    sbox_9[45] = 8'd216;
    sbox_9[46] = 8'd49;
    sbox_9[47] = 8'd21;
    sbox_9[48] = 8'd4;
    sbox_9[49] = 8'd199;
    sbox_9[50] = 8'd35;
    sbox_9[51] = 8'd195;
    sbox_9[52] = 8'd24;
    sbox_9[53] = 8'd150;
    sbox_9[54] = 8'd5;
    sbox_9[55] = 8'd154;
    sbox_9[56] = 8'd7;
    sbox_9[57] = 8'd18;
    sbox_9[58] = 8'd128;
    sbox_9[59] = 8'd226;
    sbox_9[60] = 8'd235;
    sbox_9[61] = 8'd39;
    sbox_9[62] = 8'd178;
    sbox_9[63] = 8'd117;
    sbox_9[64] = 8'd9;
    sbox_9[65] = 8'd131;
    sbox_9[66] = 8'd44;
    sbox_9[67] = 8'd26;
    sbox_9[68] = 8'd27;
    sbox_9[69] = 8'd110;
    sbox_9[70] = 8'd90;
    sbox_9[71] = 8'd160;
    sbox_9[72] = 8'd82;
    sbox_9[73] = 8'd59;
    sbox_9[74] = 8'd214;
    sbox_9[75] = 8'd179;
    sbox_9[76] = 8'd41;
    sbox_9[77] = 8'd227;
    sbox_9[78] = 8'd47;
    sbox_9[79] = 8'd132;
    sbox_9[80] = 8'd83;
    sbox_9[81] = 8'd209;
    sbox_9[82] = 8'd0;
    sbox_9[83] = 8'd237;
    sbox_9[84] = 8'd32;
    sbox_9[85] = 8'd252;
    sbox_9[86] = 8'd177;
    sbox_9[87] = 8'd91;
    sbox_9[88] = 8'd106;
    sbox_9[89] = 8'd203;
    sbox_9[90] = 8'd190;
    sbox_9[91] = 8'd57;
    sbox_9[92] = 8'd74;
    sbox_9[93] = 8'd76;
    sbox_9[94] = 8'd88;
    sbox_9[95] = 8'd207;
    sbox_9[96] = 8'd208;
    sbox_9[97] = 8'd239;
    sbox_9[98] = 8'd170;
    sbox_9[99] = 8'd251;
    sbox_9[100] = 8'd67;
    sbox_9[101] = 8'd77;
    sbox_9[102] = 8'd51;
    sbox_9[103] = 8'd133;
    sbox_9[104] = 8'd69;
    sbox_9[105] = 8'd249;
    sbox_9[106] = 8'd2;
    sbox_9[107] = 8'd127;
    sbox_9[108] = 8'd80;
    sbox_9[109] = 8'd60;
    sbox_9[110] = 8'd159;
    sbox_9[111] = 8'd168;
    sbox_9[112] = 8'd81;
    sbox_9[113] = 8'd163;
    sbox_9[114] = 8'd64;
    sbox_9[115] = 8'd143;
    sbox_9[116] = 8'd146;
    sbox_9[117] = 8'd157;
    sbox_9[118] = 8'd56;
    sbox_9[119] = 8'd245;
    sbox_9[120] = 8'd188;
    sbox_9[121] = 8'd182;
    sbox_9[122] = 8'd218;
    sbox_9[123] = 8'd33;
    sbox_9[124] = 8'd16;
    sbox_9[125] = 8'd255;
    sbox_9[126] = 8'd243;
    sbox_9[127] = 8'd210;
    sbox_9[128] = 8'd205;
    sbox_9[129] = 8'd12;
    sbox_9[130] = 8'd19;
    sbox_9[131] = 8'd236;
    sbox_9[132] = 8'd95;
    sbox_9[133] = 8'd151;
    sbox_9[134] = 8'd68;
    sbox_9[135] = 8'd23;
    sbox_9[136] = 8'd196;
    sbox_9[137] = 8'd167;
    sbox_9[138] = 8'd126;
    sbox_9[139] = 8'd61;
    sbox_9[140] = 8'd100;
    sbox_9[141] = 8'd93;
    sbox_9[142] = 8'd25;
    sbox_9[143] = 8'd115;
    sbox_9[144] = 8'd96;
    sbox_9[145] = 8'd129;
    sbox_9[146] = 8'd79;
    sbox_9[147] = 8'd220;
    sbox_9[148] = 8'd34;
    sbox_9[149] = 8'd42;
    sbox_9[150] = 8'd144;
    sbox_9[151] = 8'd136;
    sbox_9[152] = 8'd70;
    sbox_9[153] = 8'd238;
    sbox_9[154] = 8'd184;
    sbox_9[155] = 8'd20;
    sbox_9[156] = 8'd222;
    sbox_9[157] = 8'd94;
    sbox_9[158] = 8'd11;
    sbox_9[159] = 8'd219;
    sbox_9[160] = 8'd224;
    sbox_9[161] = 8'd50;
    sbox_9[162] = 8'd58;
    sbox_9[163] = 8'd10;
    sbox_9[164] = 8'd73;
    sbox_9[165] = 8'd6;
    sbox_9[166] = 8'd36;
    sbox_9[167] = 8'd92;
    sbox_9[168] = 8'd194;
    sbox_9[169] = 8'd211;
    sbox_9[170] = 8'd172;
    sbox_9[171] = 8'd98;
    sbox_9[172] = 8'd145;
    sbox_9[173] = 8'd149;
    sbox_9[174] = 8'd228;
    sbox_9[175] = 8'd121;
    sbox_9[176] = 8'd231;
    sbox_9[177] = 8'd200;
    sbox_9[178] = 8'd55;
    sbox_9[179] = 8'd109;
    sbox_9[180] = 8'd141;
    sbox_9[181] = 8'd213;
    sbox_9[182] = 8'd78;
    sbox_9[183] = 8'd169;
    sbox_9[184] = 8'd108;
    sbox_9[185] = 8'd86;
    sbox_9[186] = 8'd244;
    sbox_9[187] = 8'd234;
    sbox_9[188] = 8'd101;
    sbox_9[189] = 8'd122;
    sbox_9[190] = 8'd174;
    sbox_9[191] = 8'd8;
    sbox_9[192] = 8'd186;
    sbox_9[193] = 8'd120;
    sbox_9[194] = 8'd37;
    sbox_9[195] = 8'd46;
    sbox_9[196] = 8'd28;
    sbox_9[197] = 8'd166;
    sbox_9[198] = 8'd180;
    sbox_9[199] = 8'd198;
    sbox_9[200] = 8'd232;
    sbox_9[201] = 8'd221;
    sbox_9[202] = 8'd116;
    sbox_9[203] = 8'd31;
    sbox_9[204] = 8'd75;
    sbox_9[205] = 8'd189;
    sbox_9[206] = 8'd139;
    sbox_9[207] = 8'd138;
    sbox_9[208] = 8'd112;
    sbox_9[209] = 8'd62;
    sbox_9[210] = 8'd181;
    sbox_9[211] = 8'd102;
    sbox_9[212] = 8'd72;
    sbox_9[213] = 8'd3;
    sbox_9[214] = 8'd246;
    sbox_9[215] = 8'd14;
    sbox_9[216] = 8'd97;
    sbox_9[217] = 8'd53;
    sbox_9[218] = 8'd87;
    sbox_9[219] = 8'd185;
    sbox_9[220] = 8'd134;
    sbox_9[221] = 8'd193;
    sbox_9[222] = 8'd29;
    sbox_9[223] = 8'd158;
    sbox_9[224] = 8'd225;
    sbox_9[225] = 8'd248;
    sbox_9[226] = 8'd152;
    sbox_9[227] = 8'd17;
    sbox_9[228] = 8'd105;
    sbox_9[229] = 8'd217;
    sbox_9[230] = 8'd142;
    sbox_9[231] = 8'd148;
    sbox_9[232] = 8'd155;
    sbox_9[233] = 8'd30;
    sbox_9[234] = 8'd135;
    sbox_9[235] = 8'd233;
    sbox_9[236] = 8'd206;
    sbox_9[237] = 8'd85;
    sbox_9[238] = 8'd40;
    sbox_9[239] = 8'd223;
    sbox_9[240] = 8'd140;
    sbox_9[241] = 8'd161;
    sbox_9[242] = 8'd137;
    sbox_9[243] = 8'd13;
    sbox_9[244] = 8'd191;
    sbox_9[245] = 8'd230;
    sbox_9[246] = 8'd66;
    sbox_9[247] = 8'd104;
    sbox_9[248] = 8'd65;
    sbox_9[249] = 8'd153;
    sbox_9[250] = 8'd45;
    sbox_9[251] = 8'd15;
    sbox_9[252] = 8'd176;
    sbox_9[253] = 8'd84;
    sbox_9[254] = 8'd187;
    sbox_9[255] = 8'd22;
    sbox_10[0] = 8'd99;
    sbox_10[1] = 8'd124;
    sbox_10[2] = 8'd119;
    sbox_10[3] = 8'd123;
    sbox_10[4] = 8'd242;
    sbox_10[5] = 8'd107;
    sbox_10[6] = 8'd111;
    sbox_10[7] = 8'd197;
    sbox_10[8] = 8'd48;
    sbox_10[9] = 8'd1;
    sbox_10[10] = 8'd103;
    sbox_10[11] = 8'd43;
    sbox_10[12] = 8'd254;
    sbox_10[13] = 8'd215;
    sbox_10[14] = 8'd171;
    sbox_10[15] = 8'd118;
    sbox_10[16] = 8'd202;
    sbox_10[17] = 8'd130;
    sbox_10[18] = 8'd201;
    sbox_10[19] = 8'd125;
    sbox_10[20] = 8'd250;
    sbox_10[21] = 8'd89;
    sbox_10[22] = 8'd71;
    sbox_10[23] = 8'd240;
    sbox_10[24] = 8'd173;
    sbox_10[25] = 8'd212;
    sbox_10[26] = 8'd162;
    sbox_10[27] = 8'd175;
    sbox_10[28] = 8'd156;
    sbox_10[29] = 8'd164;
    sbox_10[30] = 8'd114;
    sbox_10[31] = 8'd192;
    sbox_10[32] = 8'd183;
    sbox_10[33] = 8'd253;
    sbox_10[34] = 8'd147;
    sbox_10[35] = 8'd38;
    sbox_10[36] = 8'd54;
    sbox_10[37] = 8'd63;
    sbox_10[38] = 8'd247;
    sbox_10[39] = 8'd204;
    sbox_10[40] = 8'd52;
    sbox_10[41] = 8'd165;
    sbox_10[42] = 8'd229;
    sbox_10[43] = 8'd241;
    sbox_10[44] = 8'd113;
    sbox_10[45] = 8'd216;
    sbox_10[46] = 8'd49;
    sbox_10[47] = 8'd21;
    sbox_10[48] = 8'd4;
    sbox_10[49] = 8'd199;
    sbox_10[50] = 8'd35;
    sbox_10[51] = 8'd195;
    sbox_10[52] = 8'd24;
    sbox_10[53] = 8'd150;
    sbox_10[54] = 8'd5;
    sbox_10[55] = 8'd154;
    sbox_10[56] = 8'd7;
    sbox_10[57] = 8'd18;
    sbox_10[58] = 8'd128;
    sbox_10[59] = 8'd226;
    sbox_10[60] = 8'd235;
    sbox_10[61] = 8'd39;
    sbox_10[62] = 8'd178;
    sbox_10[63] = 8'd117;
    sbox_10[64] = 8'd9;
    sbox_10[65] = 8'd131;
    sbox_10[66] = 8'd44;
    sbox_10[67] = 8'd26;
    sbox_10[68] = 8'd27;
    sbox_10[69] = 8'd110;
    sbox_10[70] = 8'd90;
    sbox_10[71] = 8'd160;
    sbox_10[72] = 8'd82;
    sbox_10[73] = 8'd59;
    sbox_10[74] = 8'd214;
    sbox_10[75] = 8'd179;
    sbox_10[76] = 8'd41;
    sbox_10[77] = 8'd227;
    sbox_10[78] = 8'd47;
    sbox_10[79] = 8'd132;
    sbox_10[80] = 8'd83;
    sbox_10[81] = 8'd209;
    sbox_10[82] = 8'd0;
    sbox_10[83] = 8'd237;
    sbox_10[84] = 8'd32;
    sbox_10[85] = 8'd252;
    sbox_10[86] = 8'd177;
    sbox_10[87] = 8'd91;
    sbox_10[88] = 8'd106;
    sbox_10[89] = 8'd203;
    sbox_10[90] = 8'd190;
    sbox_10[91] = 8'd57;
    sbox_10[92] = 8'd74;
    sbox_10[93] = 8'd76;
    sbox_10[94] = 8'd88;
    sbox_10[95] = 8'd207;
    sbox_10[96] = 8'd208;
    sbox_10[97] = 8'd239;
    sbox_10[98] = 8'd170;
    sbox_10[99] = 8'd251;
    sbox_10[100] = 8'd67;
    sbox_10[101] = 8'd77;
    sbox_10[102] = 8'd51;
    sbox_10[103] = 8'd133;
    sbox_10[104] = 8'd69;
    sbox_10[105] = 8'd249;
    sbox_10[106] = 8'd2;
    sbox_10[107] = 8'd127;
    sbox_10[108] = 8'd80;
    sbox_10[109] = 8'd60;
    sbox_10[110] = 8'd159;
    sbox_10[111] = 8'd168;
    sbox_10[112] = 8'd81;
    sbox_10[113] = 8'd163;
    sbox_10[114] = 8'd64;
    sbox_10[115] = 8'd143;
    sbox_10[116] = 8'd146;
    sbox_10[117] = 8'd157;
    sbox_10[118] = 8'd56;
    sbox_10[119] = 8'd245;
    sbox_10[120] = 8'd188;
    sbox_10[121] = 8'd182;
    sbox_10[122] = 8'd218;
    sbox_10[123] = 8'd33;
    sbox_10[124] = 8'd16;
    sbox_10[125] = 8'd255;
    sbox_10[126] = 8'd243;
    sbox_10[127] = 8'd210;
    sbox_10[128] = 8'd205;
    sbox_10[129] = 8'd12;
    sbox_10[130] = 8'd19;
    sbox_10[131] = 8'd236;
    sbox_10[132] = 8'd95;
    sbox_10[133] = 8'd151;
    sbox_10[134] = 8'd68;
    sbox_10[135] = 8'd23;
    sbox_10[136] = 8'd196;
    sbox_10[137] = 8'd167;
    sbox_10[138] = 8'd126;
    sbox_10[139] = 8'd61;
    sbox_10[140] = 8'd100;
    sbox_10[141] = 8'd93;
    sbox_10[142] = 8'd25;
    sbox_10[143] = 8'd115;
    sbox_10[144] = 8'd96;
    sbox_10[145] = 8'd129;
    sbox_10[146] = 8'd79;
    sbox_10[147] = 8'd220;
    sbox_10[148] = 8'd34;
    sbox_10[149] = 8'd42;
    sbox_10[150] = 8'd144;
    sbox_10[151] = 8'd136;
    sbox_10[152] = 8'd70;
    sbox_10[153] = 8'd238;
    sbox_10[154] = 8'd184;
    sbox_10[155] = 8'd20;
    sbox_10[156] = 8'd222;
    sbox_10[157] = 8'd94;
    sbox_10[158] = 8'd11;
    sbox_10[159] = 8'd219;
    sbox_10[160] = 8'd224;
    sbox_10[161] = 8'd50;
    sbox_10[162] = 8'd58;
    sbox_10[163] = 8'd10;
    sbox_10[164] = 8'd73;
    sbox_10[165] = 8'd6;
    sbox_10[166] = 8'd36;
    sbox_10[167] = 8'd92;
    sbox_10[168] = 8'd194;
    sbox_10[169] = 8'd211;
    sbox_10[170] = 8'd172;
    sbox_10[171] = 8'd98;
    sbox_10[172] = 8'd145;
    sbox_10[173] = 8'd149;
    sbox_10[174] = 8'd228;
    sbox_10[175] = 8'd121;
    sbox_10[176] = 8'd231;
    sbox_10[177] = 8'd200;
    sbox_10[178] = 8'd55;
    sbox_10[179] = 8'd109;
    sbox_10[180] = 8'd141;
    sbox_10[181] = 8'd213;
    sbox_10[182] = 8'd78;
    sbox_10[183] = 8'd169;
    sbox_10[184] = 8'd108;
    sbox_10[185] = 8'd86;
    sbox_10[186] = 8'd244;
    sbox_10[187] = 8'd234;
    sbox_10[188] = 8'd101;
    sbox_10[189] = 8'd122;
    sbox_10[190] = 8'd174;
    sbox_10[191] = 8'd8;
    sbox_10[192] = 8'd186;
    sbox_10[193] = 8'd120;
    sbox_10[194] = 8'd37;
    sbox_10[195] = 8'd46;
    sbox_10[196] = 8'd28;
    sbox_10[197] = 8'd166;
    sbox_10[198] = 8'd180;
    sbox_10[199] = 8'd198;
    sbox_10[200] = 8'd232;
    sbox_10[201] = 8'd221;
    sbox_10[202] = 8'd116;
    sbox_10[203] = 8'd31;
    sbox_10[204] = 8'd75;
    sbox_10[205] = 8'd189;
    sbox_10[206] = 8'd139;
    sbox_10[207] = 8'd138;
    sbox_10[208] = 8'd112;
    sbox_10[209] = 8'd62;
    sbox_10[210] = 8'd181;
    sbox_10[211] = 8'd102;
    sbox_10[212] = 8'd72;
    sbox_10[213] = 8'd3;
    sbox_10[214] = 8'd246;
    sbox_10[215] = 8'd14;
    sbox_10[216] = 8'd97;
    sbox_10[217] = 8'd53;
    sbox_10[218] = 8'd87;
    sbox_10[219] = 8'd185;
    sbox_10[220] = 8'd134;
    sbox_10[221] = 8'd193;
    sbox_10[222] = 8'd29;
    sbox_10[223] = 8'd158;
    sbox_10[224] = 8'd225;
    sbox_10[225] = 8'd248;
    sbox_10[226] = 8'd152;
    sbox_10[227] = 8'd17;
    sbox_10[228] = 8'd105;
    sbox_10[229] = 8'd217;
    sbox_10[230] = 8'd142;
    sbox_10[231] = 8'd148;
    sbox_10[232] = 8'd155;
    sbox_10[233] = 8'd30;
    sbox_10[234] = 8'd135;
    sbox_10[235] = 8'd233;
    sbox_10[236] = 8'd206;
    sbox_10[237] = 8'd85;
    sbox_10[238] = 8'd40;
    sbox_10[239] = 8'd223;
    sbox_10[240] = 8'd140;
    sbox_10[241] = 8'd161;
    sbox_10[242] = 8'd137;
    sbox_10[243] = 8'd13;
    sbox_10[244] = 8'd191;
    sbox_10[245] = 8'd230;
    sbox_10[246] = 8'd66;
    sbox_10[247] = 8'd104;
    sbox_10[248] = 8'd65;
    sbox_10[249] = 8'd153;
    sbox_10[250] = 8'd45;
    sbox_10[251] = 8'd15;
    sbox_10[252] = 8'd176;
    sbox_10[253] = 8'd84;
    sbox_10[254] = 8'd187;
    sbox_10[255] = 8'd22;
    sbox_11[0] = 8'd99;
    sbox_11[1] = 8'd124;
    sbox_11[2] = 8'd119;
    sbox_11[3] = 8'd123;
    sbox_11[4] = 8'd242;
    sbox_11[5] = 8'd107;
    sbox_11[6] = 8'd111;
    sbox_11[7] = 8'd197;
    sbox_11[8] = 8'd48;
    sbox_11[9] = 8'd1;
    sbox_11[10] = 8'd103;
    sbox_11[11] = 8'd43;
    sbox_11[12] = 8'd254;
    sbox_11[13] = 8'd215;
    sbox_11[14] = 8'd171;
    sbox_11[15] = 8'd118;
    sbox_11[16] = 8'd202;
    sbox_11[17] = 8'd130;
    sbox_11[18] = 8'd201;
    sbox_11[19] = 8'd125;
    sbox_11[20] = 8'd250;
    sbox_11[21] = 8'd89;
    sbox_11[22] = 8'd71;
    sbox_11[23] = 8'd240;
    sbox_11[24] = 8'd173;
    sbox_11[25] = 8'd212;
    sbox_11[26] = 8'd162;
    sbox_11[27] = 8'd175;
    sbox_11[28] = 8'd156;
    sbox_11[29] = 8'd164;
    sbox_11[30] = 8'd114;
    sbox_11[31] = 8'd192;
    sbox_11[32] = 8'd183;
    sbox_11[33] = 8'd253;
    sbox_11[34] = 8'd147;
    sbox_11[35] = 8'd38;
    sbox_11[36] = 8'd54;
    sbox_11[37] = 8'd63;
    sbox_11[38] = 8'd247;
    sbox_11[39] = 8'd204;
    sbox_11[40] = 8'd52;
    sbox_11[41] = 8'd165;
    sbox_11[42] = 8'd229;
    sbox_11[43] = 8'd241;
    sbox_11[44] = 8'd113;
    sbox_11[45] = 8'd216;
    sbox_11[46] = 8'd49;
    sbox_11[47] = 8'd21;
    sbox_11[48] = 8'd4;
    sbox_11[49] = 8'd199;
    sbox_11[50] = 8'd35;
    sbox_11[51] = 8'd195;
    sbox_11[52] = 8'd24;
    sbox_11[53] = 8'd150;
    sbox_11[54] = 8'd5;
    sbox_11[55] = 8'd154;
    sbox_11[56] = 8'd7;
    sbox_11[57] = 8'd18;
    sbox_11[58] = 8'd128;
    sbox_11[59] = 8'd226;
    sbox_11[60] = 8'd235;
    sbox_11[61] = 8'd39;
    sbox_11[62] = 8'd178;
    sbox_11[63] = 8'd117;
    sbox_11[64] = 8'd9;
    sbox_11[65] = 8'd131;
    sbox_11[66] = 8'd44;
    sbox_11[67] = 8'd26;
    sbox_11[68] = 8'd27;
    sbox_11[69] = 8'd110;
    sbox_11[70] = 8'd90;
    sbox_11[71] = 8'd160;
    sbox_11[72] = 8'd82;
    sbox_11[73] = 8'd59;
    sbox_11[74] = 8'd214;
    sbox_11[75] = 8'd179;
    sbox_11[76] = 8'd41;
    sbox_11[77] = 8'd227;
    sbox_11[78] = 8'd47;
    sbox_11[79] = 8'd132;
    sbox_11[80] = 8'd83;
    sbox_11[81] = 8'd209;
    sbox_11[82] = 8'd0;
    sbox_11[83] = 8'd237;
    sbox_11[84] = 8'd32;
    sbox_11[85] = 8'd252;
    sbox_11[86] = 8'd177;
    sbox_11[87] = 8'd91;
    sbox_11[88] = 8'd106;
    sbox_11[89] = 8'd203;
    sbox_11[90] = 8'd190;
    sbox_11[91] = 8'd57;
    sbox_11[92] = 8'd74;
    sbox_11[93] = 8'd76;
    sbox_11[94] = 8'd88;
    sbox_11[95] = 8'd207;
    sbox_11[96] = 8'd208;
    sbox_11[97] = 8'd239;
    sbox_11[98] = 8'd170;
    sbox_11[99] = 8'd251;
    sbox_11[100] = 8'd67;
    sbox_11[101] = 8'd77;
    sbox_11[102] = 8'd51;
    sbox_11[103] = 8'd133;
    sbox_11[104] = 8'd69;
    sbox_11[105] = 8'd249;
    sbox_11[106] = 8'd2;
    sbox_11[107] = 8'd127;
    sbox_11[108] = 8'd80;
    sbox_11[109] = 8'd60;
    sbox_11[110] = 8'd159;
    sbox_11[111] = 8'd168;
    sbox_11[112] = 8'd81;
    sbox_11[113] = 8'd163;
    sbox_11[114] = 8'd64;
    sbox_11[115] = 8'd143;
    sbox_11[116] = 8'd146;
    sbox_11[117] = 8'd157;
    sbox_11[118] = 8'd56;
    sbox_11[119] = 8'd245;
    sbox_11[120] = 8'd188;
    sbox_11[121] = 8'd182;
    sbox_11[122] = 8'd218;
    sbox_11[123] = 8'd33;
    sbox_11[124] = 8'd16;
    sbox_11[125] = 8'd255;
    sbox_11[126] = 8'd243;
    sbox_11[127] = 8'd210;
    sbox_11[128] = 8'd205;
    sbox_11[129] = 8'd12;
    sbox_11[130] = 8'd19;
    sbox_11[131] = 8'd236;
    sbox_11[132] = 8'd95;
    sbox_11[133] = 8'd151;
    sbox_11[134] = 8'd68;
    sbox_11[135] = 8'd23;
    sbox_11[136] = 8'd196;
    sbox_11[137] = 8'd167;
    sbox_11[138] = 8'd126;
    sbox_11[139] = 8'd61;
    sbox_11[140] = 8'd100;
    sbox_11[141] = 8'd93;
    sbox_11[142] = 8'd25;
    sbox_11[143] = 8'd115;
    sbox_11[144] = 8'd96;
    sbox_11[145] = 8'd129;
    sbox_11[146] = 8'd79;
    sbox_11[147] = 8'd220;
    sbox_11[148] = 8'd34;
    sbox_11[149] = 8'd42;
    sbox_11[150] = 8'd144;
    sbox_11[151] = 8'd136;
    sbox_11[152] = 8'd70;
    sbox_11[153] = 8'd238;
    sbox_11[154] = 8'd184;
    sbox_11[155] = 8'd20;
    sbox_11[156] = 8'd222;
    sbox_11[157] = 8'd94;
    sbox_11[158] = 8'd11;
    sbox_11[159] = 8'd219;
    sbox_11[160] = 8'd224;
    sbox_11[161] = 8'd50;
    sbox_11[162] = 8'd58;
    sbox_11[163] = 8'd10;
    sbox_11[164] = 8'd73;
    sbox_11[165] = 8'd6;
    sbox_11[166] = 8'd36;
    sbox_11[167] = 8'd92;
    sbox_11[168] = 8'd194;
    sbox_11[169] = 8'd211;
    sbox_11[170] = 8'd172;
    sbox_11[171] = 8'd98;
    sbox_11[172] = 8'd145;
    sbox_11[173] = 8'd149;
    sbox_11[174] = 8'd228;
    sbox_11[175] = 8'd121;
    sbox_11[176] = 8'd231;
    sbox_11[177] = 8'd200;
    sbox_11[178] = 8'd55;
    sbox_11[179] = 8'd109;
    sbox_11[180] = 8'd141;
    sbox_11[181] = 8'd213;
    sbox_11[182] = 8'd78;
    sbox_11[183] = 8'd169;
    sbox_11[184] = 8'd108;
    sbox_11[185] = 8'd86;
    sbox_11[186] = 8'd244;
    sbox_11[187] = 8'd234;
    sbox_11[188] = 8'd101;
    sbox_11[189] = 8'd122;
    sbox_11[190] = 8'd174;
    sbox_11[191] = 8'd8;
    sbox_11[192] = 8'd186;
    sbox_11[193] = 8'd120;
    sbox_11[194] = 8'd37;
    sbox_11[195] = 8'd46;
    sbox_11[196] = 8'd28;
    sbox_11[197] = 8'd166;
    sbox_11[198] = 8'd180;
    sbox_11[199] = 8'd198;
    sbox_11[200] = 8'd232;
    sbox_11[201] = 8'd221;
    sbox_11[202] = 8'd116;
    sbox_11[203] = 8'd31;
    sbox_11[204] = 8'd75;
    sbox_11[205] = 8'd189;
    sbox_11[206] = 8'd139;
    sbox_11[207] = 8'd138;
    sbox_11[208] = 8'd112;
    sbox_11[209] = 8'd62;
    sbox_11[210] = 8'd181;
    sbox_11[211] = 8'd102;
    sbox_11[212] = 8'd72;
    sbox_11[213] = 8'd3;
    sbox_11[214] = 8'd246;
    sbox_11[215] = 8'd14;
    sbox_11[216] = 8'd97;
    sbox_11[217] = 8'd53;
    sbox_11[218] = 8'd87;
    sbox_11[219] = 8'd185;
    sbox_11[220] = 8'd134;
    sbox_11[221] = 8'd193;
    sbox_11[222] = 8'd29;
    sbox_11[223] = 8'd158;
    sbox_11[224] = 8'd225;
    sbox_11[225] = 8'd248;
    sbox_11[226] = 8'd152;
    sbox_11[227] = 8'd17;
    sbox_11[228] = 8'd105;
    sbox_11[229] = 8'd217;
    sbox_11[230] = 8'd142;
    sbox_11[231] = 8'd148;
    sbox_11[232] = 8'd155;
    sbox_11[233] = 8'd30;
    sbox_11[234] = 8'd135;
    sbox_11[235] = 8'd233;
    sbox_11[236] = 8'd206;
    sbox_11[237] = 8'd85;
    sbox_11[238] = 8'd40;
    sbox_11[239] = 8'd223;
    sbox_11[240] = 8'd140;
    sbox_11[241] = 8'd161;
    sbox_11[242] = 8'd137;
    sbox_11[243] = 8'd13;
    sbox_11[244] = 8'd191;
    sbox_11[245] = 8'd230;
    sbox_11[246] = 8'd66;
    sbox_11[247] = 8'd104;
    sbox_11[248] = 8'd65;
    sbox_11[249] = 8'd153;
    sbox_11[250] = 8'd45;
    sbox_11[251] = 8'd15;
    sbox_11[252] = 8'd176;
    sbox_11[253] = 8'd84;
    sbox_11[254] = 8'd187;
    sbox_11[255] = 8'd22;
    sbox_12[0] = 8'd99;
    sbox_12[1] = 8'd124;
    sbox_12[2] = 8'd119;
    sbox_12[3] = 8'd123;
    sbox_12[4] = 8'd242;
    sbox_12[5] = 8'd107;
    sbox_12[6] = 8'd111;
    sbox_12[7] = 8'd197;
    sbox_12[8] = 8'd48;
    sbox_12[9] = 8'd1;
    sbox_12[10] = 8'd103;
    sbox_12[11] = 8'd43;
    sbox_12[12] = 8'd254;
    sbox_12[13] = 8'd215;
    sbox_12[14] = 8'd171;
    sbox_12[15] = 8'd118;
    sbox_12[16] = 8'd202;
    sbox_12[17] = 8'd130;
    sbox_12[18] = 8'd201;
    sbox_12[19] = 8'd125;
    sbox_12[20] = 8'd250;
    sbox_12[21] = 8'd89;
    sbox_12[22] = 8'd71;
    sbox_12[23] = 8'd240;
    sbox_12[24] = 8'd173;
    sbox_12[25] = 8'd212;
    sbox_12[26] = 8'd162;
    sbox_12[27] = 8'd175;
    sbox_12[28] = 8'd156;
    sbox_12[29] = 8'd164;
    sbox_12[30] = 8'd114;
    sbox_12[31] = 8'd192;
    sbox_12[32] = 8'd183;
    sbox_12[33] = 8'd253;
    sbox_12[34] = 8'd147;
    sbox_12[35] = 8'd38;
    sbox_12[36] = 8'd54;
    sbox_12[37] = 8'd63;
    sbox_12[38] = 8'd247;
    sbox_12[39] = 8'd204;
    sbox_12[40] = 8'd52;
    sbox_12[41] = 8'd165;
    sbox_12[42] = 8'd229;
    sbox_12[43] = 8'd241;
    sbox_12[44] = 8'd113;
    sbox_12[45] = 8'd216;
    sbox_12[46] = 8'd49;
    sbox_12[47] = 8'd21;
    sbox_12[48] = 8'd4;
    sbox_12[49] = 8'd199;
    sbox_12[50] = 8'd35;
    sbox_12[51] = 8'd195;
    sbox_12[52] = 8'd24;
    sbox_12[53] = 8'd150;
    sbox_12[54] = 8'd5;
    sbox_12[55] = 8'd154;
    sbox_12[56] = 8'd7;
    sbox_12[57] = 8'd18;
    sbox_12[58] = 8'd128;
    sbox_12[59] = 8'd226;
    sbox_12[60] = 8'd235;
    sbox_12[61] = 8'd39;
    sbox_12[62] = 8'd178;
    sbox_12[63] = 8'd117;
    sbox_12[64] = 8'd9;
    sbox_12[65] = 8'd131;
    sbox_12[66] = 8'd44;
    sbox_12[67] = 8'd26;
    sbox_12[68] = 8'd27;
    sbox_12[69] = 8'd110;
    sbox_12[70] = 8'd90;
    sbox_12[71] = 8'd160;
    sbox_12[72] = 8'd82;
    sbox_12[73] = 8'd59;
    sbox_12[74] = 8'd214;
    sbox_12[75] = 8'd179;
    sbox_12[76] = 8'd41;
    sbox_12[77] = 8'd227;
    sbox_12[78] = 8'd47;
    sbox_12[79] = 8'd132;
    sbox_12[80] = 8'd83;
    sbox_12[81] = 8'd209;
    sbox_12[82] = 8'd0;
    sbox_12[83] = 8'd237;
    sbox_12[84] = 8'd32;
    sbox_12[85] = 8'd252;
    sbox_12[86] = 8'd177;
    sbox_12[87] = 8'd91;
    sbox_12[88] = 8'd106;
    sbox_12[89] = 8'd203;
    sbox_12[90] = 8'd190;
    sbox_12[91] = 8'd57;
    sbox_12[92] = 8'd74;
    sbox_12[93] = 8'd76;
    sbox_12[94] = 8'd88;
    sbox_12[95] = 8'd207;
    sbox_12[96] = 8'd208;
    sbox_12[97] = 8'd239;
    sbox_12[98] = 8'd170;
    sbox_12[99] = 8'd251;
    sbox_12[100] = 8'd67;
    sbox_12[101] = 8'd77;
    sbox_12[102] = 8'd51;
    sbox_12[103] = 8'd133;
    sbox_12[104] = 8'd69;
    sbox_12[105] = 8'd249;
    sbox_12[106] = 8'd2;
    sbox_12[107] = 8'd127;
    sbox_12[108] = 8'd80;
    sbox_12[109] = 8'd60;
    sbox_12[110] = 8'd159;
    sbox_12[111] = 8'd168;
    sbox_12[112] = 8'd81;
    sbox_12[113] = 8'd163;
    sbox_12[114] = 8'd64;
    sbox_12[115] = 8'd143;
    sbox_12[116] = 8'd146;
    sbox_12[117] = 8'd157;
    sbox_12[118] = 8'd56;
    sbox_12[119] = 8'd245;
    sbox_12[120] = 8'd188;
    sbox_12[121] = 8'd182;
    sbox_12[122] = 8'd218;
    sbox_12[123] = 8'd33;
    sbox_12[124] = 8'd16;
    sbox_12[125] = 8'd255;
    sbox_12[126] = 8'd243;
    sbox_12[127] = 8'd210;
    sbox_12[128] = 8'd205;
    sbox_12[129] = 8'd12;
    sbox_12[130] = 8'd19;
    sbox_12[131] = 8'd236;
    sbox_12[132] = 8'd95;
    sbox_12[133] = 8'd151;
    sbox_12[134] = 8'd68;
    sbox_12[135] = 8'd23;
    sbox_12[136] = 8'd196;
    sbox_12[137] = 8'd167;
    sbox_12[138] = 8'd126;
    sbox_12[139] = 8'd61;
    sbox_12[140] = 8'd100;
    sbox_12[141] = 8'd93;
    sbox_12[142] = 8'd25;
    sbox_12[143] = 8'd115;
    sbox_12[144] = 8'd96;
    sbox_12[145] = 8'd129;
    sbox_12[146] = 8'd79;
    sbox_12[147] = 8'd220;
    sbox_12[148] = 8'd34;
    sbox_12[149] = 8'd42;
    sbox_12[150] = 8'd144;
    sbox_12[151] = 8'd136;
    sbox_12[152] = 8'd70;
    sbox_12[153] = 8'd238;
    sbox_12[154] = 8'd184;
    sbox_12[155] = 8'd20;
    sbox_12[156] = 8'd222;
    sbox_12[157] = 8'd94;
    sbox_12[158] = 8'd11;
    sbox_12[159] = 8'd219;
    sbox_12[160] = 8'd224;
    sbox_12[161] = 8'd50;
    sbox_12[162] = 8'd58;
    sbox_12[163] = 8'd10;
    sbox_12[164] = 8'd73;
    sbox_12[165] = 8'd6;
    sbox_12[166] = 8'd36;
    sbox_12[167] = 8'd92;
    sbox_12[168] = 8'd194;
    sbox_12[169] = 8'd211;
    sbox_12[170] = 8'd172;
    sbox_12[171] = 8'd98;
    sbox_12[172] = 8'd145;
    sbox_12[173] = 8'd149;
    sbox_12[174] = 8'd228;
    sbox_12[175] = 8'd121;
    sbox_12[176] = 8'd231;
    sbox_12[177] = 8'd200;
    sbox_12[178] = 8'd55;
    sbox_12[179] = 8'd109;
    sbox_12[180] = 8'd141;
    sbox_12[181] = 8'd213;
    sbox_12[182] = 8'd78;
    sbox_12[183] = 8'd169;
    sbox_12[184] = 8'd108;
    sbox_12[185] = 8'd86;
    sbox_12[186] = 8'd244;
    sbox_12[187] = 8'd234;
    sbox_12[188] = 8'd101;
    sbox_12[189] = 8'd122;
    sbox_12[190] = 8'd174;
    sbox_12[191] = 8'd8;
    sbox_12[192] = 8'd186;
    sbox_12[193] = 8'd120;
    sbox_12[194] = 8'd37;
    sbox_12[195] = 8'd46;
    sbox_12[196] = 8'd28;
    sbox_12[197] = 8'd166;
    sbox_12[198] = 8'd180;
    sbox_12[199] = 8'd198;
    sbox_12[200] = 8'd232;
    sbox_12[201] = 8'd221;
    sbox_12[202] = 8'd116;
    sbox_12[203] = 8'd31;
    sbox_12[204] = 8'd75;
    sbox_12[205] = 8'd189;
    sbox_12[206] = 8'd139;
    sbox_12[207] = 8'd138;
    sbox_12[208] = 8'd112;
    sbox_12[209] = 8'd62;
    sbox_12[210] = 8'd181;
    sbox_12[211] = 8'd102;
    sbox_12[212] = 8'd72;
    sbox_12[213] = 8'd3;
    sbox_12[214] = 8'd246;
    sbox_12[215] = 8'd14;
    sbox_12[216] = 8'd97;
    sbox_12[217] = 8'd53;
    sbox_12[218] = 8'd87;
    sbox_12[219] = 8'd185;
    sbox_12[220] = 8'd134;
    sbox_12[221] = 8'd193;
    sbox_12[222] = 8'd29;
    sbox_12[223] = 8'd158;
    sbox_12[224] = 8'd225;
    sbox_12[225] = 8'd248;
    sbox_12[226] = 8'd152;
    sbox_12[227] = 8'd17;
    sbox_12[228] = 8'd105;
    sbox_12[229] = 8'd217;
    sbox_12[230] = 8'd142;
    sbox_12[231] = 8'd148;
    sbox_12[232] = 8'd155;
    sbox_12[233] = 8'd30;
    sbox_12[234] = 8'd135;
    sbox_12[235] = 8'd233;
    sbox_12[236] = 8'd206;
    sbox_12[237] = 8'd85;
    sbox_12[238] = 8'd40;
    sbox_12[239] = 8'd223;
    sbox_12[240] = 8'd140;
    sbox_12[241] = 8'd161;
    sbox_12[242] = 8'd137;
    sbox_12[243] = 8'd13;
    sbox_12[244] = 8'd191;
    sbox_12[245] = 8'd230;
    sbox_12[246] = 8'd66;
    sbox_12[247] = 8'd104;
    sbox_12[248] = 8'd65;
    sbox_12[249] = 8'd153;
    sbox_12[250] = 8'd45;
    sbox_12[251] = 8'd15;
    sbox_12[252] = 8'd176;
    sbox_12[253] = 8'd84;
    sbox_12[254] = 8'd187;
    sbox_12[255] = 8'd22;
    sbox_13[0] = 8'd99;
    sbox_13[1] = 8'd124;
    sbox_13[2] = 8'd119;
    sbox_13[3] = 8'd123;
    sbox_13[4] = 8'd242;
    sbox_13[5] = 8'd107;
    sbox_13[6] = 8'd111;
    sbox_13[7] = 8'd197;
    sbox_13[8] = 8'd48;
    sbox_13[9] = 8'd1;
    sbox_13[10] = 8'd103;
    sbox_13[11] = 8'd43;
    sbox_13[12] = 8'd254;
    sbox_13[13] = 8'd215;
    sbox_13[14] = 8'd171;
    sbox_13[15] = 8'd118;
    sbox_13[16] = 8'd202;
    sbox_13[17] = 8'd130;
    sbox_13[18] = 8'd201;
    sbox_13[19] = 8'd125;
    sbox_13[20] = 8'd250;
    sbox_13[21] = 8'd89;
    sbox_13[22] = 8'd71;
    sbox_13[23] = 8'd240;
    sbox_13[24] = 8'd173;
    sbox_13[25] = 8'd212;
    sbox_13[26] = 8'd162;
    sbox_13[27] = 8'd175;
    sbox_13[28] = 8'd156;
    sbox_13[29] = 8'd164;
    sbox_13[30] = 8'd114;
    sbox_13[31] = 8'd192;
    sbox_13[32] = 8'd183;
    sbox_13[33] = 8'd253;
    sbox_13[34] = 8'd147;
    sbox_13[35] = 8'd38;
    sbox_13[36] = 8'd54;
    sbox_13[37] = 8'd63;
    sbox_13[38] = 8'd247;
    sbox_13[39] = 8'd204;
    sbox_13[40] = 8'd52;
    sbox_13[41] = 8'd165;
    sbox_13[42] = 8'd229;
    sbox_13[43] = 8'd241;
    sbox_13[44] = 8'd113;
    sbox_13[45] = 8'd216;
    sbox_13[46] = 8'd49;
    sbox_13[47] = 8'd21;
    sbox_13[48] = 8'd4;
    sbox_13[49] = 8'd199;
    sbox_13[50] = 8'd35;
    sbox_13[51] = 8'd195;
    sbox_13[52] = 8'd24;
    sbox_13[53] = 8'd150;
    sbox_13[54] = 8'd5;
    sbox_13[55] = 8'd154;
    sbox_13[56] = 8'd7;
    sbox_13[57] = 8'd18;
    sbox_13[58] = 8'd128;
    sbox_13[59] = 8'd226;
    sbox_13[60] = 8'd235;
    sbox_13[61] = 8'd39;
    sbox_13[62] = 8'd178;
    sbox_13[63] = 8'd117;
    sbox_13[64] = 8'd9;
    sbox_13[65] = 8'd131;
    sbox_13[66] = 8'd44;
    sbox_13[67] = 8'd26;
    sbox_13[68] = 8'd27;
    sbox_13[69] = 8'd110;
    sbox_13[70] = 8'd90;
    sbox_13[71] = 8'd160;
    sbox_13[72] = 8'd82;
    sbox_13[73] = 8'd59;
    sbox_13[74] = 8'd214;
    sbox_13[75] = 8'd179;
    sbox_13[76] = 8'd41;
    sbox_13[77] = 8'd227;
    sbox_13[78] = 8'd47;
    sbox_13[79] = 8'd132;
    sbox_13[80] = 8'd83;
    sbox_13[81] = 8'd209;
    sbox_13[82] = 8'd0;
    sbox_13[83] = 8'd237;
    sbox_13[84] = 8'd32;
    sbox_13[85] = 8'd252;
    sbox_13[86] = 8'd177;
    sbox_13[87] = 8'd91;
    sbox_13[88] = 8'd106;
    sbox_13[89] = 8'd203;
    sbox_13[90] = 8'd190;
    sbox_13[91] = 8'd57;
    sbox_13[92] = 8'd74;
    sbox_13[93] = 8'd76;
    sbox_13[94] = 8'd88;
    sbox_13[95] = 8'd207;
    sbox_13[96] = 8'd208;
    sbox_13[97] = 8'd239;
    sbox_13[98] = 8'd170;
    sbox_13[99] = 8'd251;
    sbox_13[100] = 8'd67;
    sbox_13[101] = 8'd77;
    sbox_13[102] = 8'd51;
    sbox_13[103] = 8'd133;
    sbox_13[104] = 8'd69;
    sbox_13[105] = 8'd249;
    sbox_13[106] = 8'd2;
    sbox_13[107] = 8'd127;
    sbox_13[108] = 8'd80;
    sbox_13[109] = 8'd60;
    sbox_13[110] = 8'd159;
    sbox_13[111] = 8'd168;
    sbox_13[112] = 8'd81;
    sbox_13[113] = 8'd163;
    sbox_13[114] = 8'd64;
    sbox_13[115] = 8'd143;
    sbox_13[116] = 8'd146;
    sbox_13[117] = 8'd157;
    sbox_13[118] = 8'd56;
    sbox_13[119] = 8'd245;
    sbox_13[120] = 8'd188;
    sbox_13[121] = 8'd182;
    sbox_13[122] = 8'd218;
    sbox_13[123] = 8'd33;
    sbox_13[124] = 8'd16;
    sbox_13[125] = 8'd255;
    sbox_13[126] = 8'd243;
    sbox_13[127] = 8'd210;
    sbox_13[128] = 8'd205;
    sbox_13[129] = 8'd12;
    sbox_13[130] = 8'd19;
    sbox_13[131] = 8'd236;
    sbox_13[132] = 8'd95;
    sbox_13[133] = 8'd151;
    sbox_13[134] = 8'd68;
    sbox_13[135] = 8'd23;
    sbox_13[136] = 8'd196;
    sbox_13[137] = 8'd167;
    sbox_13[138] = 8'd126;
    sbox_13[139] = 8'd61;
    sbox_13[140] = 8'd100;
    sbox_13[141] = 8'd93;
    sbox_13[142] = 8'd25;
    sbox_13[143] = 8'd115;
    sbox_13[144] = 8'd96;
    sbox_13[145] = 8'd129;
    sbox_13[146] = 8'd79;
    sbox_13[147] = 8'd220;
    sbox_13[148] = 8'd34;
    sbox_13[149] = 8'd42;
    sbox_13[150] = 8'd144;
    sbox_13[151] = 8'd136;
    sbox_13[152] = 8'd70;
    sbox_13[153] = 8'd238;
    sbox_13[154] = 8'd184;
    sbox_13[155] = 8'd20;
    sbox_13[156] = 8'd222;
    sbox_13[157] = 8'd94;
    sbox_13[158] = 8'd11;
    sbox_13[159] = 8'd219;
    sbox_13[160] = 8'd224;
    sbox_13[161] = 8'd50;
    sbox_13[162] = 8'd58;
    sbox_13[163] = 8'd10;
    sbox_13[164] = 8'd73;
    sbox_13[165] = 8'd6;
    sbox_13[166] = 8'd36;
    sbox_13[167] = 8'd92;
    sbox_13[168] = 8'd194;
    sbox_13[169] = 8'd211;
    sbox_13[170] = 8'd172;
    sbox_13[171] = 8'd98;
    sbox_13[172] = 8'd145;
    sbox_13[173] = 8'd149;
    sbox_13[174] = 8'd228;
    sbox_13[175] = 8'd121;
    sbox_13[176] = 8'd231;
    sbox_13[177] = 8'd200;
    sbox_13[178] = 8'd55;
    sbox_13[179] = 8'd109;
    sbox_13[180] = 8'd141;
    sbox_13[181] = 8'd213;
    sbox_13[182] = 8'd78;
    sbox_13[183] = 8'd169;
    sbox_13[184] = 8'd108;
    sbox_13[185] = 8'd86;
    sbox_13[186] = 8'd244;
    sbox_13[187] = 8'd234;
    sbox_13[188] = 8'd101;
    sbox_13[189] = 8'd122;
    sbox_13[190] = 8'd174;
    sbox_13[191] = 8'd8;
    sbox_13[192] = 8'd186;
    sbox_13[193] = 8'd120;
    sbox_13[194] = 8'd37;
    sbox_13[195] = 8'd46;
    sbox_13[196] = 8'd28;
    sbox_13[197] = 8'd166;
    sbox_13[198] = 8'd180;
    sbox_13[199] = 8'd198;
    sbox_13[200] = 8'd232;
    sbox_13[201] = 8'd221;
    sbox_13[202] = 8'd116;
    sbox_13[203] = 8'd31;
    sbox_13[204] = 8'd75;
    sbox_13[205] = 8'd189;
    sbox_13[206] = 8'd139;
    sbox_13[207] = 8'd138;
    sbox_13[208] = 8'd112;
    sbox_13[209] = 8'd62;
    sbox_13[210] = 8'd181;
    sbox_13[211] = 8'd102;
    sbox_13[212] = 8'd72;
    sbox_13[213] = 8'd3;
    sbox_13[214] = 8'd246;
    sbox_13[215] = 8'd14;
    sbox_13[216] = 8'd97;
    sbox_13[217] = 8'd53;
    sbox_13[218] = 8'd87;
    sbox_13[219] = 8'd185;
    sbox_13[220] = 8'd134;
    sbox_13[221] = 8'd193;
    sbox_13[222] = 8'd29;
    sbox_13[223] = 8'd158;
    sbox_13[224] = 8'd225;
    sbox_13[225] = 8'd248;
    sbox_13[226] = 8'd152;
    sbox_13[227] = 8'd17;
    sbox_13[228] = 8'd105;
    sbox_13[229] = 8'd217;
    sbox_13[230] = 8'd142;
    sbox_13[231] = 8'd148;
    sbox_13[232] = 8'd155;
    sbox_13[233] = 8'd30;
    sbox_13[234] = 8'd135;
    sbox_13[235] = 8'd233;
    sbox_13[236] = 8'd206;
    sbox_13[237] = 8'd85;
    sbox_13[238] = 8'd40;
    sbox_13[239] = 8'd223;
    sbox_13[240] = 8'd140;
    sbox_13[241] = 8'd161;
    sbox_13[242] = 8'd137;
    sbox_13[243] = 8'd13;
    sbox_13[244] = 8'd191;
    sbox_13[245] = 8'd230;
    sbox_13[246] = 8'd66;
    sbox_13[247] = 8'd104;
    sbox_13[248] = 8'd65;
    sbox_13[249] = 8'd153;
    sbox_13[250] = 8'd45;
    sbox_13[251] = 8'd15;
    sbox_13[252] = 8'd176;
    sbox_13[253] = 8'd84;
    sbox_13[254] = 8'd187;
    sbox_13[255] = 8'd22;
    sbox_14[0] = 8'd99;
    sbox_14[1] = 8'd124;
    sbox_14[2] = 8'd119;
    sbox_14[3] = 8'd123;
    sbox_14[4] = 8'd242;
    sbox_14[5] = 8'd107;
    sbox_14[6] = 8'd111;
    sbox_14[7] = 8'd197;
    sbox_14[8] = 8'd48;
    sbox_14[9] = 8'd1;
    sbox_14[10] = 8'd103;
    sbox_14[11] = 8'd43;
    sbox_14[12] = 8'd254;
    sbox_14[13] = 8'd215;
    sbox_14[14] = 8'd171;
    sbox_14[15] = 8'd118;
    sbox_14[16] = 8'd202;
    sbox_14[17] = 8'd130;
    sbox_14[18] = 8'd201;
    sbox_14[19] = 8'd125;
    sbox_14[20] = 8'd250;
    sbox_14[21] = 8'd89;
    sbox_14[22] = 8'd71;
    sbox_14[23] = 8'd240;
    sbox_14[24] = 8'd173;
    sbox_14[25] = 8'd212;
    sbox_14[26] = 8'd162;
    sbox_14[27] = 8'd175;
    sbox_14[28] = 8'd156;
    sbox_14[29] = 8'd164;
    sbox_14[30] = 8'd114;
    sbox_14[31] = 8'd192;
    sbox_14[32] = 8'd183;
    sbox_14[33] = 8'd253;
    sbox_14[34] = 8'd147;
    sbox_14[35] = 8'd38;
    sbox_14[36] = 8'd54;
    sbox_14[37] = 8'd63;
    sbox_14[38] = 8'd247;
    sbox_14[39] = 8'd204;
    sbox_14[40] = 8'd52;
    sbox_14[41] = 8'd165;
    sbox_14[42] = 8'd229;
    sbox_14[43] = 8'd241;
    sbox_14[44] = 8'd113;
    sbox_14[45] = 8'd216;
    sbox_14[46] = 8'd49;
    sbox_14[47] = 8'd21;
    sbox_14[48] = 8'd4;
    sbox_14[49] = 8'd199;
    sbox_14[50] = 8'd35;
    sbox_14[51] = 8'd195;
    sbox_14[52] = 8'd24;
    sbox_14[53] = 8'd150;
    sbox_14[54] = 8'd5;
    sbox_14[55] = 8'd154;
    sbox_14[56] = 8'd7;
    sbox_14[57] = 8'd18;
    sbox_14[58] = 8'd128;
    sbox_14[59] = 8'd226;
    sbox_14[60] = 8'd235;
    sbox_14[61] = 8'd39;
    sbox_14[62] = 8'd178;
    sbox_14[63] = 8'd117;
    sbox_14[64] = 8'd9;
    sbox_14[65] = 8'd131;
    sbox_14[66] = 8'd44;
    sbox_14[67] = 8'd26;
    sbox_14[68] = 8'd27;
    sbox_14[69] = 8'd110;
    sbox_14[70] = 8'd90;
    sbox_14[71] = 8'd160;
    sbox_14[72] = 8'd82;
    sbox_14[73] = 8'd59;
    sbox_14[74] = 8'd214;
    sbox_14[75] = 8'd179;
    sbox_14[76] = 8'd41;
    sbox_14[77] = 8'd227;
    sbox_14[78] = 8'd47;
    sbox_14[79] = 8'd132;
    sbox_14[80] = 8'd83;
    sbox_14[81] = 8'd209;
    sbox_14[82] = 8'd0;
    sbox_14[83] = 8'd237;
    sbox_14[84] = 8'd32;
    sbox_14[85] = 8'd252;
    sbox_14[86] = 8'd177;
    sbox_14[87] = 8'd91;
    sbox_14[88] = 8'd106;
    sbox_14[89] = 8'd203;
    sbox_14[90] = 8'd190;
    sbox_14[91] = 8'd57;
    sbox_14[92] = 8'd74;
    sbox_14[93] = 8'd76;
    sbox_14[94] = 8'd88;
    sbox_14[95] = 8'd207;
    sbox_14[96] = 8'd208;
    sbox_14[97] = 8'd239;
    sbox_14[98] = 8'd170;
    sbox_14[99] = 8'd251;
    sbox_14[100] = 8'd67;
    sbox_14[101] = 8'd77;
    sbox_14[102] = 8'd51;
    sbox_14[103] = 8'd133;
    sbox_14[104] = 8'd69;
    sbox_14[105] = 8'd249;
    sbox_14[106] = 8'd2;
    sbox_14[107] = 8'd127;
    sbox_14[108] = 8'd80;
    sbox_14[109] = 8'd60;
    sbox_14[110] = 8'd159;
    sbox_14[111] = 8'd168;
    sbox_14[112] = 8'd81;
    sbox_14[113] = 8'd163;
    sbox_14[114] = 8'd64;
    sbox_14[115] = 8'd143;
    sbox_14[116] = 8'd146;
    sbox_14[117] = 8'd157;
    sbox_14[118] = 8'd56;
    sbox_14[119] = 8'd245;
    sbox_14[120] = 8'd188;
    sbox_14[121] = 8'd182;
    sbox_14[122] = 8'd218;
    sbox_14[123] = 8'd33;
    sbox_14[124] = 8'd16;
    sbox_14[125] = 8'd255;
    sbox_14[126] = 8'd243;
    sbox_14[127] = 8'd210;
    sbox_14[128] = 8'd205;
    sbox_14[129] = 8'd12;
    sbox_14[130] = 8'd19;
    sbox_14[131] = 8'd236;
    sbox_14[132] = 8'd95;
    sbox_14[133] = 8'd151;
    sbox_14[134] = 8'd68;
    sbox_14[135] = 8'd23;
    sbox_14[136] = 8'd196;
    sbox_14[137] = 8'd167;
    sbox_14[138] = 8'd126;
    sbox_14[139] = 8'd61;
    sbox_14[140] = 8'd100;
    sbox_14[141] = 8'd93;
    sbox_14[142] = 8'd25;
    sbox_14[143] = 8'd115;
    sbox_14[144] = 8'd96;
    sbox_14[145] = 8'd129;
    sbox_14[146] = 8'd79;
    sbox_14[147] = 8'd220;
    sbox_14[148] = 8'd34;
    sbox_14[149] = 8'd42;
    sbox_14[150] = 8'd144;
    sbox_14[151] = 8'd136;
    sbox_14[152] = 8'd70;
    sbox_14[153] = 8'd238;
    sbox_14[154] = 8'd184;
    sbox_14[155] = 8'd20;
    sbox_14[156] = 8'd222;
    sbox_14[157] = 8'd94;
    sbox_14[158] = 8'd11;
    sbox_14[159] = 8'd219;
    sbox_14[160] = 8'd224;
    sbox_14[161] = 8'd50;
    sbox_14[162] = 8'd58;
    sbox_14[163] = 8'd10;
    sbox_14[164] = 8'd73;
    sbox_14[165] = 8'd6;
    sbox_14[166] = 8'd36;
    sbox_14[167] = 8'd92;
    sbox_14[168] = 8'd194;
    sbox_14[169] = 8'd211;
    sbox_14[170] = 8'd172;
    sbox_14[171] = 8'd98;
    sbox_14[172] = 8'd145;
    sbox_14[173] = 8'd149;
    sbox_14[174] = 8'd228;
    sbox_14[175] = 8'd121;
    sbox_14[176] = 8'd231;
    sbox_14[177] = 8'd200;
    sbox_14[178] = 8'd55;
    sbox_14[179] = 8'd109;
    sbox_14[180] = 8'd141;
    sbox_14[181] = 8'd213;
    sbox_14[182] = 8'd78;
    sbox_14[183] = 8'd169;
    sbox_14[184] = 8'd108;
    sbox_14[185] = 8'd86;
    sbox_14[186] = 8'd244;
    sbox_14[187] = 8'd234;
    sbox_14[188] = 8'd101;
    sbox_14[189] = 8'd122;
    sbox_14[190] = 8'd174;
    sbox_14[191] = 8'd8;
    sbox_14[192] = 8'd186;
    sbox_14[193] = 8'd120;
    sbox_14[194] = 8'd37;
    sbox_14[195] = 8'd46;
    sbox_14[196] = 8'd28;
    sbox_14[197] = 8'd166;
    sbox_14[198] = 8'd180;
    sbox_14[199] = 8'd198;
    sbox_14[200] = 8'd232;
    sbox_14[201] = 8'd221;
    sbox_14[202] = 8'd116;
    sbox_14[203] = 8'd31;
    sbox_14[204] = 8'd75;
    sbox_14[205] = 8'd189;
    sbox_14[206] = 8'd139;
    sbox_14[207] = 8'd138;
    sbox_14[208] = 8'd112;
    sbox_14[209] = 8'd62;
    sbox_14[210] = 8'd181;
    sbox_14[211] = 8'd102;
    sbox_14[212] = 8'd72;
    sbox_14[213] = 8'd3;
    sbox_14[214] = 8'd246;
    sbox_14[215] = 8'd14;
    sbox_14[216] = 8'd97;
    sbox_14[217] = 8'd53;
    sbox_14[218] = 8'd87;
    sbox_14[219] = 8'd185;
    sbox_14[220] = 8'd134;
    sbox_14[221] = 8'd193;
    sbox_14[222] = 8'd29;
    sbox_14[223] = 8'd158;
    sbox_14[224] = 8'd225;
    sbox_14[225] = 8'd248;
    sbox_14[226] = 8'd152;
    sbox_14[227] = 8'd17;
    sbox_14[228] = 8'd105;
    sbox_14[229] = 8'd217;
    sbox_14[230] = 8'd142;
    sbox_14[231] = 8'd148;
    sbox_14[232] = 8'd155;
    sbox_14[233] = 8'd30;
    sbox_14[234] = 8'd135;
    sbox_14[235] = 8'd233;
    sbox_14[236] = 8'd206;
    sbox_14[237] = 8'd85;
    sbox_14[238] = 8'd40;
    sbox_14[239] = 8'd223;
    sbox_14[240] = 8'd140;
    sbox_14[241] = 8'd161;
    sbox_14[242] = 8'd137;
    sbox_14[243] = 8'd13;
    sbox_14[244] = 8'd191;
    sbox_14[245] = 8'd230;
    sbox_14[246] = 8'd66;
    sbox_14[247] = 8'd104;
    sbox_14[248] = 8'd65;
    sbox_14[249] = 8'd153;
    sbox_14[250] = 8'd45;
    sbox_14[251] = 8'd15;
    sbox_14[252] = 8'd176;
    sbox_14[253] = 8'd84;
    sbox_14[254] = 8'd187;
    sbox_14[255] = 8'd22;
    sbox_15[0] = 8'd99;
    sbox_15[1] = 8'd124;
    sbox_15[2] = 8'd119;
    sbox_15[3] = 8'd123;
    sbox_15[4] = 8'd242;
    sbox_15[5] = 8'd107;
    sbox_15[6] = 8'd111;
    sbox_15[7] = 8'd197;
    sbox_15[8] = 8'd48;
    sbox_15[9] = 8'd1;
    sbox_15[10] = 8'd103;
    sbox_15[11] = 8'd43;
    sbox_15[12] = 8'd254;
    sbox_15[13] = 8'd215;
    sbox_15[14] = 8'd171;
    sbox_15[15] = 8'd118;
    sbox_15[16] = 8'd202;
    sbox_15[17] = 8'd130;
    sbox_15[18] = 8'd201;
    sbox_15[19] = 8'd125;
    sbox_15[20] = 8'd250;
    sbox_15[21] = 8'd89;
    sbox_15[22] = 8'd71;
    sbox_15[23] = 8'd240;
    sbox_15[24] = 8'd173;
    sbox_15[25] = 8'd212;
    sbox_15[26] = 8'd162;
    sbox_15[27] = 8'd175;
    sbox_15[28] = 8'd156;
    sbox_15[29] = 8'd164;
    sbox_15[30] = 8'd114;
    sbox_15[31] = 8'd192;
    sbox_15[32] = 8'd183;
    sbox_15[33] = 8'd253;
    sbox_15[34] = 8'd147;
    sbox_15[35] = 8'd38;
    sbox_15[36] = 8'd54;
    sbox_15[37] = 8'd63;
    sbox_15[38] = 8'd247;
    sbox_15[39] = 8'd204;
    sbox_15[40] = 8'd52;
    sbox_15[41] = 8'd165;
    sbox_15[42] = 8'd229;
    sbox_15[43] = 8'd241;
    sbox_15[44] = 8'd113;
    sbox_15[45] = 8'd216;
    sbox_15[46] = 8'd49;
    sbox_15[47] = 8'd21;
    sbox_15[48] = 8'd4;
    sbox_15[49] = 8'd199;
    sbox_15[50] = 8'd35;
    sbox_15[51] = 8'd195;
    sbox_15[52] = 8'd24;
    sbox_15[53] = 8'd150;
    sbox_15[54] = 8'd5;
    sbox_15[55] = 8'd154;
    sbox_15[56] = 8'd7;
    sbox_15[57] = 8'd18;
    sbox_15[58] = 8'd128;
    sbox_15[59] = 8'd226;
    sbox_15[60] = 8'd235;
    sbox_15[61] = 8'd39;
    sbox_15[62] = 8'd178;
    sbox_15[63] = 8'd117;
    sbox_15[64] = 8'd9;
    sbox_15[65] = 8'd131;
    sbox_15[66] = 8'd44;
    sbox_15[67] = 8'd26;
    sbox_15[68] = 8'd27;
    sbox_15[69] = 8'd110;
    sbox_15[70] = 8'd90;
    sbox_15[71] = 8'd160;
    sbox_15[72] = 8'd82;
    sbox_15[73] = 8'd59;
    sbox_15[74] = 8'd214;
    sbox_15[75] = 8'd179;
    sbox_15[76] = 8'd41;
    sbox_15[77] = 8'd227;
    sbox_15[78] = 8'd47;
    sbox_15[79] = 8'd132;
    sbox_15[80] = 8'd83;
    sbox_15[81] = 8'd209;
    sbox_15[82] = 8'd0;
    sbox_15[83] = 8'd237;
    sbox_15[84] = 8'd32;
    sbox_15[85] = 8'd252;
    sbox_15[86] = 8'd177;
    sbox_15[87] = 8'd91;
    sbox_15[88] = 8'd106;
    sbox_15[89] = 8'd203;
    sbox_15[90] = 8'd190;
    sbox_15[91] = 8'd57;
    sbox_15[92] = 8'd74;
    sbox_15[93] = 8'd76;
    sbox_15[94] = 8'd88;
    sbox_15[95] = 8'd207;
    sbox_15[96] = 8'd208;
    sbox_15[97] = 8'd239;
    sbox_15[98] = 8'd170;
    sbox_15[99] = 8'd251;
    sbox_15[100] = 8'd67;
    sbox_15[101] = 8'd77;
    sbox_15[102] = 8'd51;
    sbox_15[103] = 8'd133;
    sbox_15[104] = 8'd69;
    sbox_15[105] = 8'd249;
    sbox_15[106] = 8'd2;
    sbox_15[107] = 8'd127;
    sbox_15[108] = 8'd80;
    sbox_15[109] = 8'd60;
    sbox_15[110] = 8'd159;
    sbox_15[111] = 8'd168;
    sbox_15[112] = 8'd81;
    sbox_15[113] = 8'd163;
    sbox_15[114] = 8'd64;
    sbox_15[115] = 8'd143;
    sbox_15[116] = 8'd146;
    sbox_15[117] = 8'd157;
    sbox_15[118] = 8'd56;
    sbox_15[119] = 8'd245;
    sbox_15[120] = 8'd188;
    sbox_15[121] = 8'd182;
    sbox_15[122] = 8'd218;
    sbox_15[123] = 8'd33;
    sbox_15[124] = 8'd16;
    sbox_15[125] = 8'd255;
    sbox_15[126] = 8'd243;
    sbox_15[127] = 8'd210;
    sbox_15[128] = 8'd205;
    sbox_15[129] = 8'd12;
    sbox_15[130] = 8'd19;
    sbox_15[131] = 8'd236;
    sbox_15[132] = 8'd95;
    sbox_15[133] = 8'd151;
    sbox_15[134] = 8'd68;
    sbox_15[135] = 8'd23;
    sbox_15[136] = 8'd196;
    sbox_15[137] = 8'd167;
    sbox_15[138] = 8'd126;
    sbox_15[139] = 8'd61;
    sbox_15[140] = 8'd100;
    sbox_15[141] = 8'd93;
    sbox_15[142] = 8'd25;
    sbox_15[143] = 8'd115;
    sbox_15[144] = 8'd96;
    sbox_15[145] = 8'd129;
    sbox_15[146] = 8'd79;
    sbox_15[147] = 8'd220;
    sbox_15[148] = 8'd34;
    sbox_15[149] = 8'd42;
    sbox_15[150] = 8'd144;
    sbox_15[151] = 8'd136;
    sbox_15[152] = 8'd70;
    sbox_15[153] = 8'd238;
    sbox_15[154] = 8'd184;
    sbox_15[155] = 8'd20;
    sbox_15[156] = 8'd222;
    sbox_15[157] = 8'd94;
    sbox_15[158] = 8'd11;
    sbox_15[159] = 8'd219;
    sbox_15[160] = 8'd224;
    sbox_15[161] = 8'd50;
    sbox_15[162] = 8'd58;
    sbox_15[163] = 8'd10;
    sbox_15[164] = 8'd73;
    sbox_15[165] = 8'd6;
    sbox_15[166] = 8'd36;
    sbox_15[167] = 8'd92;
    sbox_15[168] = 8'd194;
    sbox_15[169] = 8'd211;
    sbox_15[170] = 8'd172;
    sbox_15[171] = 8'd98;
    sbox_15[172] = 8'd145;
    sbox_15[173] = 8'd149;
    sbox_15[174] = 8'd228;
    sbox_15[175] = 8'd121;
    sbox_15[176] = 8'd231;
    sbox_15[177] = 8'd200;
    sbox_15[178] = 8'd55;
    sbox_15[179] = 8'd109;
    sbox_15[180] = 8'd141;
    sbox_15[181] = 8'd213;
    sbox_15[182] = 8'd78;
    sbox_15[183] = 8'd169;
    sbox_15[184] = 8'd108;
    sbox_15[185] = 8'd86;
    sbox_15[186] = 8'd244;
    sbox_15[187] = 8'd234;
    sbox_15[188] = 8'd101;
    sbox_15[189] = 8'd122;
    sbox_15[190] = 8'd174;
    sbox_15[191] = 8'd8;
    sbox_15[192] = 8'd186;
    sbox_15[193] = 8'd120;
    sbox_15[194] = 8'd37;
    sbox_15[195] = 8'd46;
    sbox_15[196] = 8'd28;
    sbox_15[197] = 8'd166;
    sbox_15[198] = 8'd180;
    sbox_15[199] = 8'd198;
    sbox_15[200] = 8'd232;
    sbox_15[201] = 8'd221;
    sbox_15[202] = 8'd116;
    sbox_15[203] = 8'd31;
    sbox_15[204] = 8'd75;
    sbox_15[205] = 8'd189;
    sbox_15[206] = 8'd139;
    sbox_15[207] = 8'd138;
    sbox_15[208] = 8'd112;
    sbox_15[209] = 8'd62;
    sbox_15[210] = 8'd181;
    sbox_15[211] = 8'd102;
    sbox_15[212] = 8'd72;
    sbox_15[213] = 8'd3;
    sbox_15[214] = 8'd246;
    sbox_15[215] = 8'd14;
    sbox_15[216] = 8'd97;
    sbox_15[217] = 8'd53;
    sbox_15[218] = 8'd87;
    sbox_15[219] = 8'd185;
    sbox_15[220] = 8'd134;
    sbox_15[221] = 8'd193;
    sbox_15[222] = 8'd29;
    sbox_15[223] = 8'd158;
    sbox_15[224] = 8'd225;
    sbox_15[225] = 8'd248;
    sbox_15[226] = 8'd152;
    sbox_15[227] = 8'd17;
    sbox_15[228] = 8'd105;
    sbox_15[229] = 8'd217;
    sbox_15[230] = 8'd142;
    sbox_15[231] = 8'd148;
    sbox_15[232] = 8'd155;
    sbox_15[233] = 8'd30;
    sbox_15[234] = 8'd135;
    sbox_15[235] = 8'd233;
    sbox_15[236] = 8'd206;
    sbox_15[237] = 8'd85;
    sbox_15[238] = 8'd40;
    sbox_15[239] = 8'd223;
    sbox_15[240] = 8'd140;
    sbox_15[241] = 8'd161;
    sbox_15[242] = 8'd137;
    sbox_15[243] = 8'd13;
    sbox_15[244] = 8'd191;
    sbox_15[245] = 8'd230;
    sbox_15[246] = 8'd66;
    sbox_15[247] = 8'd104;
    sbox_15[248] = 8'd65;
    sbox_15[249] = 8'd153;
    sbox_15[250] = 8'd45;
    sbox_15[251] = 8'd15;
    sbox_15[252] = 8'd176;
    sbox_15[253] = 8'd84;
    sbox_15[254] = 8'd187;
    sbox_15[255] = 8'd22;
end
    assign lookup_sbox_0_enable = ((control_274_0)||((control_274_1)||((control_274_5)||((control_274_6)||((control_274_10)||((control_274_11)||((control_274_16)||((control_274_19)||((control_274_17)||((control_274_21)||((control_274_22)||((control_274_28)||((control_274_26)||((control_274_27)||((control_274_37)||((control_274_32)||((control_274_38)||((control_274_46)||((control_274_44)||((control_274_43)||((control_274_55)||((control_274_48)||((control_274_49)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))))))))))))))))))));
    assign lookup_sbox_0_0 = ((control_274_0)?({(operation_274_124[111:104])}):((control_274_1)?({(operation_274_119[7:0])}):((control_274_5)?({(operation_274_1821[7:0])}):((control_274_6)?({(operation_274_1749[7:0])}):((control_274_10)?({(operation_274_1699[7:0])}):((control_274_11)?({(operation_274_2250[7:0])}):((control_274_16)?({(operation_274_2679[7:0])}):((control_274_19)?({(operation_274_2128[7:0])}):((control_274_17)?({(operation_274_2607[7:0])}):((control_274_21)?({(operation_274_3108[7:0])}):((control_274_22)?({(operation_274_3109[7:0])}):((control_274_28)?({(operation_274_2557[7:0])}):((control_274_26)?({(operation_274_3537[7:0])}):((control_274_27)?({(operation_274_3538[7:0])}):((control_274_37)?({(operation_274_2986[7:0])}):((control_274_32)?({(operation_274_3966[7:0])}):((control_274_38)?({(operation_274_4395[7:0])}):((control_274_46)?({(operation_274_3415[7:0])}):((control_274_44)?({(operation_274_4752[7:0])}):((control_274_43)?({(operation_274_4824[7:0])}):((control_274_55)?({(operation_274_3844[7:0])}):((control_274_48)?({(operation_274_5253[7:0])}):((control_274_49)?({(operation_274_5254[7:0])}):((control_274_64)?({(operation_274_4273[7:0])}):((control_274_73)?({(operation_274_4702[7:0])}):((control_274_82)?({(operation_274_5131[7:0])}):(1'd0)))))))))))))))))))))))))));
    assign lookup_sbox_1_enable = ((control_274_0)||((control_274_1)||((control_274_5)||((control_274_10)||((control_274_11)||((control_274_19)||((control_274_16)||((control_274_22)||((control_274_21)||((control_274_28)||((control_274_27)||((control_274_37)||((control_274_32)||((control_274_38)||((control_274_46)||((control_274_43)||((control_274_55)||((control_274_48)||((control_274_49)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))))))))))))))));
    assign lookup_sbox_1_0 = ((control_274_0)?({(operation_274_124[127:120])}):((control_274_1)?({(operation_274_103[7:0])}):((control_274_5)?({(operation_274_1822[7:0])}):((control_274_10)?({(operation_274_1700[7:0])}):((control_274_11)?({(operation_274_2232[7:0])}):((control_274_19)?({(operation_274_2129[7:0])}):((control_274_16)?({(operation_274_2680[7:0])}):((control_274_22)?({(operation_274_3036[7:0])}):((control_274_21)?({(operation_274_3090[7:0])}):((control_274_28)?({(operation_274_2558[7:0])}):((control_274_27)?({(operation_274_3519[7:0])}):((control_274_37)?({(operation_274_2987[7:0])}):((control_274_32)?({(operation_274_3948[7:0])}):((control_274_38)?({(operation_274_4396[7:0])}):((control_274_46)?({(operation_274_3416[7:0])}):((control_274_43)?({(operation_274_4806[7:0])}):((control_274_55)?({(operation_274_3845[7:0])}):((control_274_48)?({(operation_274_5235[7:0])}):((control_274_49)?({(operation_274_5181[7:0])}):((control_274_64)?({(operation_274_4274[7:0])}):((control_274_73)?({(operation_274_4703[7:0])}):((control_274_82)?({(operation_274_5132[7:0])}):(1'd0)))))))))))))))))))))));
    assign lookup_sbox_2_enable = ((control_274_0)||((control_274_1)||((control_274_5)||((control_274_10)||((control_274_11)||((control_274_19)||((control_274_16)||((control_274_28)||((control_274_27)||((control_274_37)||((control_274_32)||((control_274_38)||((control_274_46)||((control_274_43)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))))))))))));
    assign lookup_sbox_2_0 = ((control_274_0)?({(operation_274_124[119:112])}):((control_274_1)?({(operation_274_87[7:0])}):((control_274_5)?({(operation_274_1803[7:0])}):((control_274_10)?({(operation_274_1701[7:0])}):((control_274_11)?({(operation_274_2251[7:0])}):((control_274_19)?({(operation_274_2130[7:0])}):((control_274_16)?({(operation_274_2661[7:0])}):((control_274_28)?({(operation_274_2559[7:0])}):((control_274_27)?({(operation_274_3465[7:0])}):((control_274_37)?({(operation_274_2988[7:0])}):((control_274_32)?({(operation_274_3967[7:0])}):((control_274_38)?({(operation_274_4377[7:0])}):((control_274_46)?({(operation_274_3417[7:0])}):((control_274_43)?({(operation_274_4825[7:0])}):((control_274_55)?({(operation_274_3846[7:0])}):((control_274_64)?({(operation_274_4275[7:0])}):((control_274_73)?({(operation_274_4704[7:0])}):((control_274_82)?({(operation_274_5133[7:0])}):(1'd0)))))))))))))))))));
    assign lookup_sbox_3_enable = ((control_274_0)||((control_274_1)||((control_274_10)||((control_274_11)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_32)||((control_274_38)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))))))));
    assign lookup_sbox_3_0 = ((control_274_0)?({(operation_274_124[103:96])}):((control_274_1)?({(operation_274_71[7:0])}):((control_274_10)?({(operation_274_1702[7:0])}):((control_274_11)?({(operation_274_2178[7:0])}):((control_274_19)?({(operation_274_2131[7:0])}):((control_274_28)?({(operation_274_2560[7:0])}):((control_274_37)?({(operation_274_2989[7:0])}):((control_274_32)?({(operation_274_3894[7:0])}):((control_274_38)?({(operation_274_4323[7:0])}):((control_274_46)?({(operation_274_3418[7:0])}):((control_274_55)?({(operation_274_3847[7:0])}):((control_274_64)?({(operation_274_4276[7:0])}):((control_274_73)?({(operation_274_4705[7:0])}):((control_274_82)?({(operation_274_5134[7:0])}):(1'd0)))))))))))))));
    assign lookup_sbox_4_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_4_0 = ((control_274_1)?({(operation_274_55[7:0])}):((control_274_10)?({(operation_274_1703[7:0])}):((control_274_19)?({(operation_274_2132[7:0])}):((control_274_28)?({(operation_274_2561[7:0])}):((control_274_37)?({(operation_274_2990[7:0])}):((control_274_46)?({(operation_274_3419[7:0])}):((control_274_55)?({(operation_274_3848[7:0])}):((control_274_64)?({(operation_274_4277[7:0])}):((control_274_73)?({(operation_274_4706[7:0])}):((control_274_82)?({(operation_274_5135[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_5_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_5_0 = ((control_274_1)?({(operation_274_39[7:0])}):((control_274_10)?({(operation_274_1704[7:0])}):((control_274_19)?({(operation_274_2133[7:0])}):((control_274_28)?({(operation_274_2562[7:0])}):((control_274_37)?({(operation_274_2991[7:0])}):((control_274_46)?({(operation_274_3420[7:0])}):((control_274_55)?({(operation_274_3849[7:0])}):((control_274_64)?({(operation_274_4278[7:0])}):((control_274_73)?({(operation_274_4707[7:0])}):((control_274_82)?({(operation_274_5136[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_6_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_6_0 = ((control_274_1)?({(operation_274_23[7:0])}):((control_274_10)?({(operation_274_1705[7:0])}):((control_274_19)?({(operation_274_2134[7:0])}):((control_274_28)?({(operation_274_2563[7:0])}):((control_274_37)?({(operation_274_2992[7:0])}):((control_274_46)?({(operation_274_3421[7:0])}):((control_274_55)?({(operation_274_3850[7:0])}):((control_274_64)?({(operation_274_4279[7:0])}):((control_274_73)?({(operation_274_4708[7:0])}):((control_274_82)?({(operation_274_5137[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_7_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_7_0 = ((control_274_1)?({(operation_274_7[7:0])}):((control_274_10)?({(operation_274_1706[7:0])}):((control_274_19)?({(operation_274_2135[7:0])}):((control_274_28)?({(operation_274_2564[7:0])}):((control_274_37)?({(operation_274_2993[7:0])}):((control_274_46)?({(operation_274_3422[7:0])}):((control_274_55)?({(operation_274_3851[7:0])}):((control_274_64)?({(operation_274_4280[7:0])}):((control_274_73)?({(operation_274_4709[7:0])}):((control_274_82)?({(operation_274_5138[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_8_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_8_0 = ((control_274_1)?({(operation_274_15[7:0])}):((control_274_10)?({(operation_274_1707[7:0])}):((control_274_19)?({(operation_274_2136[7:0])}):((control_274_28)?({(operation_274_2565[7:0])}):((control_274_37)?({(operation_274_2994[7:0])}):((control_274_46)?({(operation_274_3423[7:0])}):((control_274_55)?({(operation_274_3852[7:0])}):((control_274_64)?({(operation_274_4281[7:0])}):((control_274_73)?({(operation_274_4710[7:0])}):((control_274_82)?({(operation_274_5139[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_9_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_9_0 = ((control_274_1)?({(operation_274_31[7:0])}):((control_274_10)?({(operation_274_1708[7:0])}):((control_274_19)?({(operation_274_2137[7:0])}):((control_274_28)?({(operation_274_2566[7:0])}):((control_274_37)?({(operation_274_2995[7:0])}):((control_274_46)?({(operation_274_3424[7:0])}):((control_274_55)?({(operation_274_3853[7:0])}):((control_274_64)?({(operation_274_4282[7:0])}):((control_274_73)?({(operation_274_4711[7:0])}):((control_274_82)?({(operation_274_5140[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_10_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_10_0 = ((control_274_1)?({(operation_274_47[7:0])}):((control_274_10)?({(operation_274_1709[7:0])}):((control_274_19)?({(operation_274_2138[7:0])}):((control_274_28)?({(operation_274_2567[7:0])}):((control_274_37)?({(operation_274_2996[7:0])}):((control_274_46)?({(operation_274_3425[7:0])}):((control_274_55)?({(operation_274_3854[7:0])}):((control_274_64)?({(operation_274_4283[7:0])}):((control_274_73)?({(operation_274_4712[7:0])}):((control_274_82)?({(operation_274_5141[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_11_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_11_0 = ((control_274_1)?({(operation_274_63[7:0])}):((control_274_10)?({(operation_274_1710[7:0])}):((control_274_19)?({(operation_274_2139[7:0])}):((control_274_28)?({(operation_274_2568[7:0])}):((control_274_37)?({(operation_274_2997[7:0])}):((control_274_46)?({(operation_274_3426[7:0])}):((control_274_55)?({(operation_274_3855[7:0])}):((control_274_64)?({(operation_274_4284[7:0])}):((control_274_73)?({(operation_274_4713[7:0])}):((control_274_82)?({(operation_274_5142[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_12_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_12_0 = ((control_274_1)?({(operation_274_79[7:0])}):((control_274_10)?({(operation_274_1711[7:0])}):((control_274_19)?({(operation_274_2140[7:0])}):((control_274_28)?({(operation_274_2569[7:0])}):((control_274_37)?({(operation_274_2998[7:0])}):((control_274_46)?({(operation_274_3427[7:0])}):((control_274_55)?({(operation_274_3856[7:0])}):((control_274_64)?({(operation_274_4285[7:0])}):((control_274_73)?({(operation_274_4714[7:0])}):((control_274_82)?({(operation_274_5143[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_13_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_13_0 = ((control_274_1)?({(operation_274_95[7:0])}):((control_274_10)?({(operation_274_1712[7:0])}):((control_274_19)?({(operation_274_2141[7:0])}):((control_274_28)?({(operation_274_2570[7:0])}):((control_274_37)?({(operation_274_2999[7:0])}):((control_274_46)?({(operation_274_3428[7:0])}):((control_274_55)?({(operation_274_3857[7:0])}):((control_274_64)?({(operation_274_4286[7:0])}):((control_274_73)?({(operation_274_4715[7:0])}):((control_274_82)?({(operation_274_5144[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_14_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_14_0 = ((control_274_1)?({(operation_274_111[7:0])}):((control_274_10)?({(operation_274_1713[7:0])}):((control_274_19)?({(operation_274_2142[7:0])}):((control_274_28)?({(operation_274_2571[7:0])}):((control_274_37)?({(operation_274_3000[7:0])}):((control_274_46)?({(operation_274_3429[7:0])}):((control_274_55)?({(operation_274_3858[7:0])}):((control_274_64)?({(operation_274_4287[7:0])}):((control_274_73)?({(operation_274_4716[7:0])}):((control_274_82)?({(operation_274_5145[7:0])}):(1'd0)))))))))));
    assign lookup_sbox_15_enable = ((control_274_1)||((control_274_10)||((control_274_19)||((control_274_28)||((control_274_37)||((control_274_46)||((control_274_55)||((control_274_64)||((control_274_73)||((control_274_82)||(1'd0)))))))))));
    assign lookup_sbox_15_0 = ((control_274_1)?({(operation_274_127[7:0])}):((control_274_10)?({(operation_274_1714[7:0])}):((control_274_19)?({(operation_274_2143[7:0])}):((control_274_28)?({(operation_274_2572[7:0])}):((control_274_37)?({(operation_274_3001[7:0])}):((control_274_46)?({(operation_274_3430[7:0])}):((control_274_55)?({(operation_274_3859[7:0])}):((control_274_64)?({(operation_274_4288[7:0])}):((control_274_73)?({(operation_274_4717[7:0])}):((control_274_82)?({(operation_274_5146[7:0])}):(1'd0)))))))))));
    assign input_key_274 = ((start)?(key):(input_key_274_follow));
    assign input_in_274 = ((start)?(in):(input_in_274_follow));
    assign return_274 = ({(operation_274_1689[7:0]),(operation_274_1681[7:0]),(operation_274_1673[7:0]),(operation_274_1665[7:0]),(operation_274_1657[7:0]),(operation_274_1649[7:0]),(operation_274_1641[7:0]),(operation_274_1633[7:0]),(operation_274_1625[7:0]),(operation_274_1617[7:0]),(operation_274_1609[7:0]),(operation_274_1601[7:0]),(operation_274_1593[7:0]),(operation_274_1585[7:0]),(operation_274_1577[7:0]),(operation_274_1569[7:0])});
    assign operation_274_1665 = (operation_274_1664);
    assign operation_274_1689 = (operation_274_1688);
    assign operation_274_1673 = (operation_274_1672);
    assign operation_274_1633 = (operation_274_1632);
    assign operation_274_1681 = (operation_274_1680);
    assign operation_274_1657 = (operation_274_1656);
    assign operation_274_1641 = (operation_274_1640);
    assign operation_274_1601 = (operation_274_1600);
    assign operation_274_1649 = (operation_274_1648);
    assign operation_274_1625 = (operation_274_1624);
    assign operation_274_1609 = (operation_274_1608);
    assign operation_274_1569 = (operation_274_1568);
    assign operation_274_1617 = (operation_274_1616);
    assign operation_274_1593 = (operation_274_1592);
    assign operation_274_1577 = (operation_274_1576);
    assign operation_274_1585 = (operation_274_1584);
    assign operation_274_1685 = ({(operation_274_1323[7:0])});
    assign operation_274_1669 = ({(operation_274_1273[7:0])});
    assign operation_274_1653 = ({(operation_274_1303[7:0])});
    assign operation_274_1637 = ({(operation_274_1333[7:0])});
    assign operation_274_1621 = ({(operation_274_1283[7:0])});
    assign operation_274_1605 = ({(operation_274_1313[7:0])});
    assign operation_274_1589 = ({(operation_274_1343[7:0])});
    assign operation_274_1573 = ({(operation_274_1293[7:0])});
    assign operation_274_1565 = ({(operation_274_1268[7:0])});
    assign operation_274_1581 = ({(operation_274_1318[7:0])});
    assign operation_274_1597 = ({(operation_274_1288[7:0])});
    assign operation_274_1613 = ({(operation_274_1338[7:0])});
    assign operation_274_1629 = ({(operation_274_1308[7:0])});
    assign operation_274_1645 = ({(operation_274_1278[7:0])});
    assign operation_274_1661 = ({(operation_274_1328[7:0])});
    assign operation_274_1677 = ({(operation_274_1298[7:0])});
    assign operation_274_1338 = ((control_274_83)?(lookup_sbox_0_output):(operation_274_1338_latch));
    assign operation_274_1328 = ((control_274_83)?(lookup_sbox_1_output):(operation_274_1328_latch));
    assign operation_274_1318 = ((control_274_83)?(lookup_sbox_2_output):(operation_274_1318_latch));
    assign operation_274_1308 = ((control_274_83)?(lookup_sbox_3_output):(operation_274_1308_latch));
    assign operation_274_1298 = ((control_274_83)?(lookup_sbox_4_output):(operation_274_1298_latch));
    assign operation_274_1288 = ((control_274_83)?(lookup_sbox_5_output):(operation_274_1288_latch));
    assign operation_274_1278 = ((control_274_83)?(lookup_sbox_6_output):(operation_274_1278_latch));
    assign operation_274_1268 = ((control_274_83)?(lookup_sbox_7_output):(operation_274_1268_latch));
    assign operation_274_1273 = ((control_274_83)?(lookup_sbox_8_output):(operation_274_1273_latch));
    assign operation_274_1283 = ((control_274_83)?(lookup_sbox_9_output):(operation_274_1283_latch));
    assign operation_274_1293 = ((control_274_83)?(lookup_sbox_10_output):(operation_274_1293_latch));
    assign operation_274_1303 = ((control_274_83)?(lookup_sbox_11_output):(operation_274_1303_latch));
    assign operation_274_1313 = ((control_274_83)?(lookup_sbox_12_output):(operation_274_1313_latch));
    assign operation_274_1323 = ((control_274_83)?(lookup_sbox_13_output):(operation_274_1323_latch));
    assign operation_274_1333 = ((control_274_83)?(lookup_sbox_14_output):(operation_274_1333_latch));
    assign operation_274_1343 = ((control_274_83)?(lookup_sbox_15_output):(operation_274_1343_latch));
    assign operation_274_5146 = (operation_274_5162);
    assign operation_274_5145 = (operation_274_5161);
    assign operation_274_5144 = (operation_274_5160);
    assign operation_274_5143 = (operation_274_5159);
    assign operation_274_5142 = (operation_274_5158);
    assign operation_274_5141 = (operation_274_5157);
    assign operation_274_5140 = (operation_274_5156);
    assign operation_274_5139 = (operation_274_5155);
    assign operation_274_5138 = (operation_274_5154);
    assign operation_274_5137 = (operation_274_5153);
    assign operation_274_5136 = (operation_274_5152);
    assign operation_274_5135 = (operation_274_5151);
    assign operation_274_5134 = (operation_274_5150);
    assign operation_274_5133 = (operation_274_5149);
    assign operation_274_5132 = (operation_274_5148);
    assign operation_274_5131 = (operation_274_5147);
    assign operation_274_5180 = ({(operation_274_5182[7:0])});
    assign operation_274_5179 = ({(operation_274_5183[7:0])});
    assign operation_274_5178 = ({(operation_274_5184[7:0])});
    assign operation_274_5177 = ({(operation_274_5185[7:0])});
    assign operation_274_5176 = ({(operation_274_5186[7:0])});
    assign operation_274_5175 = ({(operation_274_5187[7:0])});
    assign operation_274_5174 = ({(operation_274_5188[7:0])});
    assign operation_274_5173 = ({(operation_274_5189[7:0])});
    assign operation_274_5171 = ({(operation_274_5190[7:0])});
    assign operation_274_5170 = ({(operation_274_5191[7:0])});
    assign operation_274_5169 = ({(operation_274_5192[7:0])});
    assign operation_274_5168 = ({(operation_274_5193[7:0])});
    assign operation_274_5167 = ({(operation_274_5194[7:0])});
    assign operation_274_5166 = ({(operation_274_5195[7:0])});
    assign operation_274_5165 = ({(operation_274_5196[7:0])});
    assign operation_274_5163 = ({(operation_274_5197[7:0])});
    assign operation_274_5197 = (operation_274_5214);
    assign operation_274_5196 = (operation_274_5213);
    assign operation_274_5195 = (operation_274_5212);
    assign operation_274_5194 = (operation_274_5211);
    assign operation_274_5193 = (operation_274_5210);
    assign operation_274_5192 = (operation_274_5209);
    assign operation_274_5191 = (operation_274_5208);
    assign operation_274_5190 = (operation_274_5207);
    assign operation_274_5189 = (operation_274_5206);
    assign operation_274_5188 = (operation_274_5205);
    assign operation_274_5187 = (operation_274_5204);
    assign operation_274_5186 = (operation_274_5203);
    assign operation_274_5185 = (operation_274_5202);
    assign operation_274_5184 = (operation_274_5201);
    assign operation_274_5183 = (operation_274_5200);
    assign operation_274_5182 = (operation_274_5199);
    assign operation_274_5232 = ({(operation_274_5252[7:0])});
    assign operation_274_5231 = ({(operation_274_5251[7:0])});
    assign operation_274_5230 = ({(operation_274_5250[7:0])});
    assign operation_274_5229 = ({(operation_274_5249[7:0])});
    assign operation_274_5228 = ({(operation_274_5248[7:0])});
    assign operation_274_5227 = ({(operation_274_5247[7:0])});
    assign operation_274_5226 = ({(operation_274_5246[7:0])});
    assign operation_274_5225 = ({(operation_274_5245[7:0])});
    assign operation_274_5224 = ({(operation_274_5244[7:0])});
    assign operation_274_5223 = ({(operation_274_5243[7:0])});
    assign operation_274_5222 = ({(operation_274_5242[7:0])});
    assign operation_274_5221 = ({(operation_274_5241[7:0])});
    assign operation_274_5220 = ({(operation_274_5240[7:0])});
    assign operation_274_5219 = ({(operation_274_5239[7:0])});
    assign operation_274_5218 = ({(operation_274_5238[7:0])});
    assign operation_274_5217 = ({(operation_274_5237[7:0])});
    assign operation_274_5252 = (operation_274_5272);
    assign operation_274_5251 = (operation_274_5271);
    assign operation_274_5250 = (operation_274_5270);
    assign operation_274_5249 = (operation_274_5269);
    assign operation_274_5248 = (operation_274_5268);
    assign operation_274_5247 = (operation_274_5267);
    assign operation_274_5246 = (operation_274_5266);
    assign operation_274_5245 = (operation_274_5265);
    assign operation_274_5244 = (operation_274_5264);
    assign operation_274_5243 = (operation_274_5263);
    assign operation_274_5242 = (operation_274_5262);
    assign operation_274_5241 = (operation_274_5261);
    assign operation_274_5240 = (operation_274_5260);
    assign operation_274_5239 = (operation_274_5259);
    assign operation_274_5238 = (operation_274_5258);
    assign operation_274_5237 = (operation_274_5257);
    assign operation_274_5292 = ({(operation_274_5312[7:0])});
    assign operation_274_5291 = ({(operation_274_5311[7:0])});
    assign operation_274_5290 = ({(operation_274_5310[7:0])});
    assign operation_274_5289 = ({(operation_274_5309[7:0])});
    assign operation_274_5288 = ({(operation_274_5308[7:0])});
    assign operation_274_5287 = ({(operation_274_5307[7:0])});
    assign operation_274_5286 = ({(operation_274_5306[7:0])});
    assign operation_274_5285 = ({(operation_274_5305[7:0])});
    assign operation_274_5284 = ({(operation_274_5304[7:0])});
    assign operation_274_5283 = ({(operation_274_5303[7:0])});
    assign operation_274_5282 = ({(operation_274_5302[7:0])});
    assign operation_274_5281 = ({(operation_274_5301[7:0])});
    assign operation_274_5280 = ({(operation_274_5300[7:0])});
    assign operation_274_5279 = ({(operation_274_5299[7:0])});
    assign operation_274_5278 = ({(operation_274_5298[7:0])});
    assign operation_274_5277 = ({(operation_274_5297[7:0])});
    assign operation_274_5312 = (operation_274_5332);
    assign operation_274_5311 = (operation_274_5331);
    assign operation_274_5310 = (operation_274_5330);
    assign operation_274_5309 = (operation_274_5329);
    assign operation_274_5308 = (operation_274_5328);
    assign operation_274_5307 = (operation_274_5327);
    assign operation_274_5306 = (operation_274_5326);
    assign operation_274_5305 = (operation_274_5325);
    assign operation_274_5304 = (operation_274_5324);
    assign operation_274_5303 = (operation_274_5323);
    assign operation_274_5302 = (operation_274_5322);
    assign operation_274_5301 = (operation_274_5321);
    assign operation_274_5300 = (operation_274_5320);
    assign operation_274_5299 = (operation_274_5319);
    assign operation_274_5298 = (operation_274_5318);
    assign operation_274_5297 = (operation_274_5317);
    assign operation_274_5360 = ({(operation_274_5415[7:0])});
    assign operation_274_5359 = ({(operation_274_5382[7:0])});
    assign operation_274_5358 = ({(operation_274_5416[7:0])});
    assign operation_274_5357 = ({(operation_274_5381[7:0])});
    assign operation_274_5416 = (operation_274_5440);
    assign operation_274_5415 = (operation_274_5439);
    assign operation_274_5382 = (operation_274_5422);
    assign operation_274_5381 = (operation_274_5421);
    assign operation_274_5438 = ({(operation_274_5462[7:0])});
    assign operation_274_5437 = ({(operation_274_5461[7:0])});
    assign operation_274_5436 = ({(operation_274_5460[7:0])});
    assign operation_274_5435 = ({(operation_274_5459[7:0])});
    assign operation_274_5434 = ({(operation_274_5458[7:0])});
    assign operation_274_5433 = ({(operation_274_5457[7:0])});
    assign operation_274_5432 = ({(operation_274_5456[7:0])});
    assign operation_274_5431 = ({(operation_274_5455[7:0])});
    assign operation_274_5430 = ({(operation_274_5454[7:0])});
    assign operation_274_5429 = ({(operation_274_5453[7:0])});
    assign operation_274_5428 = ({(operation_274_5452[7:0])});
    assign operation_274_5427 = ({(operation_274_5451[7:0])});
    assign operation_274_5426 = ({(operation_274_5450[7:0])});
    assign operation_274_5425 = ({(operation_274_5449[7:0])});
    assign operation_274_5424 = ({(operation_274_5448[7:0])});
    assign operation_274_5423 = ({(operation_274_5447[7:0])});
    assign operation_274_5462 = (operation_274_5485);
    assign operation_274_5461 = (operation_274_5470);
    assign operation_274_5460 = (operation_274_5484);
    assign operation_274_5459 = (operation_274_5483);
    assign operation_274_5458 = (operation_274_5482);
    assign operation_274_5457 = (operation_274_5471);
    assign operation_274_5456 = (operation_274_5481);
    assign operation_274_5455 = (operation_274_5480);
    assign operation_274_5454 = (operation_274_5479);
    assign operation_274_5453 = (operation_274_5478);
    assign operation_274_5452 = (operation_274_5477);
    assign operation_274_5451 = (operation_274_5476);
    assign operation_274_5450 = (operation_274_5475);
    assign operation_274_5449 = (operation_274_5474);
    assign operation_274_5448 = (operation_274_5473);
    assign operation_274_5447 = (operation_274_5472);
    assign operation_274_5507 = ({(operation_274_5534[7:0])});
    assign operation_274_5506 = ({(operation_274_5529[7:0])});
    assign operation_274_5505 = ({(operation_274_5530[7:0])});
    assign operation_274_5504 = ({(operation_274_5533[7:0])});
    assign operation_274_5503 = ({(operation_274_5536[7:0])});
    assign operation_274_5502 = ({(operation_274_5531[7:0])});
    assign operation_274_5501 = ({(operation_274_5532[7:0])});
    assign operation_274_5500 = ({(operation_274_5535[7:0])});
    assign operation_274_5499 = ({(operation_274_5526[7:0])});
    assign operation_274_5498 = ({(operation_274_5521[7:0])});
    assign operation_274_5497 = ({(operation_274_5524[7:0])});
    assign operation_274_5496 = ({(operation_274_5527[7:0])});
    assign operation_274_5495 = ({(operation_274_5522[7:0])});
    assign operation_274_5494 = ({(operation_274_5525[7:0])});
    assign operation_274_5493 = ({(operation_274_5528[7:0])});
    assign operation_274_5492 = ({(operation_274_5523[7:0])});
    assign operation_274_5536 = ((control_274_74)?(lookup_sbox_0_output):(operation_274_5536_latch));
    assign operation_274_5535 = ((control_274_74)?(lookup_sbox_1_output):(operation_274_5535_latch));
    assign operation_274_5534 = ((control_274_74)?(lookup_sbox_2_output):(operation_274_5534_latch));
    assign operation_274_5533 = ((control_274_74)?(lookup_sbox_3_output):(operation_274_5533_latch));
    assign operation_274_5532 = ((control_274_74)?(lookup_sbox_4_output):(operation_274_5532_latch));
    assign operation_274_5531 = ((control_274_74)?(lookup_sbox_5_output):(operation_274_5531_latch));
    assign operation_274_5530 = ((control_274_74)?(lookup_sbox_6_output):(operation_274_5530_latch));
    assign operation_274_5529 = ((control_274_74)?(lookup_sbox_7_output):(operation_274_5529_latch));
    assign operation_274_5528 = ((control_274_74)?(lookup_sbox_8_output):(operation_274_5528_latch));
    assign operation_274_5527 = ((control_274_74)?(lookup_sbox_9_output):(operation_274_5527_latch));
    assign operation_274_5526 = ((control_274_74)?(lookup_sbox_10_output):(operation_274_5526_latch));
    assign operation_274_5525 = ((control_274_74)?(lookup_sbox_11_output):(operation_274_5525_latch));
    assign operation_274_5524 = ((control_274_74)?(lookup_sbox_12_output):(operation_274_5524_latch));
    assign operation_274_5523 = ((control_274_74)?(lookup_sbox_13_output):(operation_274_5523_latch));
    assign operation_274_5522 = ((control_274_74)?(lookup_sbox_14_output):(operation_274_5522_latch));
    assign operation_274_5521 = ((control_274_74)?(lookup_sbox_15_output):(operation_274_5521_latch));
    assign operation_274_4717 = (operation_274_4733);
    assign operation_274_4716 = (operation_274_4732);
    assign operation_274_4715 = (operation_274_4731);
    assign operation_274_4714 = (operation_274_4730);
    assign operation_274_4713 = (operation_274_4729);
    assign operation_274_4712 = (operation_274_4728);
    assign operation_274_4711 = (operation_274_4727);
    assign operation_274_4710 = (operation_274_4726);
    assign operation_274_4709 = (operation_274_4725);
    assign operation_274_4708 = (operation_274_4724);
    assign operation_274_4707 = (operation_274_4723);
    assign operation_274_4706 = (operation_274_4722);
    assign operation_274_4705 = (operation_274_4721);
    assign operation_274_4704 = (operation_274_4720);
    assign operation_274_4703 = (operation_274_4719);
    assign operation_274_4702 = (operation_274_4718);
    assign operation_274_4751 = ({(operation_274_4753[7:0])});
    assign operation_274_4750 = ({(operation_274_4754[7:0])});
    assign operation_274_4749 = ({(operation_274_4755[7:0])});
    assign operation_274_4748 = ({(operation_274_4756[7:0])});
    assign operation_274_4747 = ({(operation_274_4757[7:0])});
    assign operation_274_4746 = ({(operation_274_4758[7:0])});
    assign operation_274_4745 = ({(operation_274_4759[7:0])});
    assign operation_274_4744 = ({(operation_274_4760[7:0])});
    assign operation_274_4742 = ({(operation_274_4761[7:0])});
    assign operation_274_4741 = ({(operation_274_4762[7:0])});
    assign operation_274_4740 = ({(operation_274_4763[7:0])});
    assign operation_274_4739 = ({(operation_274_4764[7:0])});
    assign operation_274_4738 = ({(operation_274_4765[7:0])});
    assign operation_274_4737 = ({(operation_274_4766[7:0])});
    assign operation_274_4736 = ({(operation_274_4767[7:0])});
    assign operation_274_4734 = ({(operation_274_4768[7:0])});
    assign operation_274_4768 = (operation_274_4785);
    assign operation_274_4767 = (operation_274_4784);
    assign operation_274_4766 = (operation_274_4783);
    assign operation_274_4765 = (operation_274_4782);
    assign operation_274_4764 = (operation_274_4781);
    assign operation_274_4763 = (operation_274_4780);
    assign operation_274_4762 = (operation_274_4779);
    assign operation_274_4761 = (operation_274_4778);
    assign operation_274_4760 = (operation_274_4777);
    assign operation_274_4759 = (operation_274_4776);
    assign operation_274_4758 = (operation_274_4775);
    assign operation_274_4757 = (operation_274_4774);
    assign operation_274_4756 = (operation_274_4773);
    assign operation_274_4755 = (operation_274_4772);
    assign operation_274_4754 = (operation_274_4771);
    assign operation_274_4753 = (operation_274_4770);
    assign operation_274_4803 = ({(operation_274_4823[7:0])});
    assign operation_274_4802 = ({(operation_274_4822[7:0])});
    assign operation_274_4801 = ({(operation_274_4821[7:0])});
    assign operation_274_4800 = ({(operation_274_4820[7:0])});
    assign operation_274_4799 = ({(operation_274_4819[7:0])});
    assign operation_274_4798 = ({(operation_274_4818[7:0])});
    assign operation_274_4797 = ({(operation_274_4817[7:0])});
    assign operation_274_4796 = ({(operation_274_4816[7:0])});
    assign operation_274_4795 = ({(operation_274_4815[7:0])});
    assign operation_274_4794 = ({(operation_274_4814[7:0])});
    assign operation_274_4793 = ({(operation_274_4813[7:0])});
    assign operation_274_4792 = ({(operation_274_4812[7:0])});
    assign operation_274_4791 = ({(operation_274_4811[7:0])});
    assign operation_274_4790 = ({(operation_274_4810[7:0])});
    assign operation_274_4789 = ({(operation_274_4809[7:0])});
    assign operation_274_4788 = ({(operation_274_4808[7:0])});
    assign operation_274_4823 = (operation_274_4843);
    assign operation_274_4822 = (operation_274_4842);
    assign operation_274_4821 = (operation_274_4841);
    assign operation_274_4820 = (operation_274_4840);
    assign operation_274_4819 = (operation_274_4839);
    assign operation_274_4818 = (operation_274_4838);
    assign operation_274_4817 = (operation_274_4837);
    assign operation_274_4816 = (operation_274_4836);
    assign operation_274_4815 = (operation_274_4835);
    assign operation_274_4814 = (operation_274_4834);
    assign operation_274_4813 = (operation_274_4833);
    assign operation_274_4812 = (operation_274_4832);
    assign operation_274_4811 = (operation_274_4831);
    assign operation_274_4810 = (operation_274_4830);
    assign operation_274_4809 = (operation_274_4829);
    assign operation_274_4808 = (operation_274_4828);
    assign operation_274_4863 = ({(operation_274_4883[7:0])});
    assign operation_274_4862 = ({(operation_274_4882[7:0])});
    assign operation_274_4861 = ({(operation_274_4881[7:0])});
    assign operation_274_4860 = ({(operation_274_4880[7:0])});
    assign operation_274_4859 = ({(operation_274_4879[7:0])});
    assign operation_274_4858 = ({(operation_274_4878[7:0])});
    assign operation_274_4857 = ({(operation_274_4877[7:0])});
    assign operation_274_4856 = ({(operation_274_4876[7:0])});
    assign operation_274_4855 = ({(operation_274_4875[7:0])});
    assign operation_274_4854 = ({(operation_274_4874[7:0])});
    assign operation_274_4853 = ({(operation_274_4873[7:0])});
    assign operation_274_4852 = ({(operation_274_4872[7:0])});
    assign operation_274_4851 = ({(operation_274_4871[7:0])});
    assign operation_274_4850 = ({(operation_274_4870[7:0])});
    assign operation_274_4849 = ({(operation_274_4869[7:0])});
    assign operation_274_4848 = ({(operation_274_4868[7:0])});
    assign operation_274_4883 = (operation_274_4903);
    assign operation_274_4882 = (operation_274_4902);
    assign operation_274_4881 = (operation_274_4901);
    assign operation_274_4880 = (operation_274_4900);
    assign operation_274_4879 = (operation_274_4899);
    assign operation_274_4878 = (operation_274_4898);
    assign operation_274_4877 = (operation_274_4897);
    assign operation_274_4876 = (operation_274_4896);
    assign operation_274_4875 = (operation_274_4895);
    assign operation_274_4874 = (operation_274_4894);
    assign operation_274_4873 = (operation_274_4893);
    assign operation_274_4872 = (operation_274_4892);
    assign operation_274_4871 = (operation_274_4891);
    assign operation_274_4870 = (operation_274_4890);
    assign operation_274_4869 = (operation_274_4889);
    assign operation_274_4868 = (operation_274_4888);
    assign operation_274_4931 = ({(operation_274_4986[7:0])});
    assign operation_274_4930 = ({(operation_274_4953[7:0])});
    assign operation_274_4929 = ({(operation_274_4987[7:0])});
    assign operation_274_4928 = ({(operation_274_4952[7:0])});
    assign operation_274_4987 = (operation_274_5011);
    assign operation_274_4986 = (operation_274_5010);
    assign operation_274_4953 = (operation_274_4993);
    assign operation_274_4952 = (operation_274_4992);
    assign operation_274_5009 = ({(operation_274_5033[7:0])});
    assign operation_274_5008 = ({(operation_274_5032[7:0])});
    assign operation_274_5007 = ({(operation_274_5031[7:0])});
    assign operation_274_5006 = ({(operation_274_5030[7:0])});
    assign operation_274_5005 = ({(operation_274_5029[7:0])});
    assign operation_274_5004 = ({(operation_274_5028[7:0])});
    assign operation_274_5003 = ({(operation_274_5027[7:0])});
    assign operation_274_5002 = ({(operation_274_5026[7:0])});
    assign operation_274_5001 = ({(operation_274_5025[7:0])});
    assign operation_274_5000 = ({(operation_274_5024[7:0])});
    assign operation_274_4999 = ({(operation_274_5023[7:0])});
    assign operation_274_4998 = ({(operation_274_5022[7:0])});
    assign operation_274_4997 = ({(operation_274_5021[7:0])});
    assign operation_274_4996 = ({(operation_274_5020[7:0])});
    assign operation_274_4995 = ({(operation_274_5019[7:0])});
    assign operation_274_4994 = ({(operation_274_5018[7:0])});
    assign operation_274_5033 = (operation_274_5056);
    assign operation_274_5032 = (operation_274_5041);
    assign operation_274_5031 = (operation_274_5055);
    assign operation_274_5030 = (operation_274_5054);
    assign operation_274_5029 = (operation_274_5053);
    assign operation_274_5028 = (operation_274_5042);
    assign operation_274_5027 = (operation_274_5052);
    assign operation_274_5026 = (operation_274_5051);
    assign operation_274_5025 = (operation_274_5050);
    assign operation_274_5024 = (operation_274_5049);
    assign operation_274_5023 = (operation_274_5048);
    assign operation_274_5022 = (operation_274_5047);
    assign operation_274_5021 = (operation_274_5046);
    assign operation_274_5020 = (operation_274_5045);
    assign operation_274_5019 = (operation_274_5044);
    assign operation_274_5018 = (operation_274_5043);
    assign operation_274_1663 = ({(operation_274_1537[7:0])});
    assign operation_274_1687 = ({(operation_274_1561[7:0])});
    assign operation_274_1537 = (operation_274_1536);
    assign operation_274_1561 = (operation_274_1560);
    assign operation_274_5078 = ({(operation_274_5105[7:0])});
    assign operation_274_5077 = ({(operation_274_5100[7:0])});
    assign operation_274_5076 = ({(operation_274_5101[7:0])});
    assign operation_274_5075 = ({(operation_274_5104[7:0])});
    assign operation_274_5074 = ({(operation_274_5107[7:0])});
    assign operation_274_5073 = ({(operation_274_5102[7:0])});
    assign operation_274_5072 = ({(operation_274_5103[7:0])});
    assign operation_274_5071 = ({(operation_274_5106[7:0])});
    assign operation_274_5070 = ({(operation_274_5097[7:0])});
    assign operation_274_5069 = ({(operation_274_5092[7:0])});
    assign operation_274_5068 = ({(operation_274_5095[7:0])});
    assign operation_274_5067 = ({(operation_274_5098[7:0])});
    assign operation_274_5066 = ({(operation_274_5093[7:0])});
    assign operation_274_5065 = ({(operation_274_5096[7:0])});
    assign operation_274_5064 = ({(operation_274_5099[7:0])});
    assign operation_274_5063 = ({(operation_274_5094[7:0])});
    assign operation_274_5107 = ((control_274_65)?(lookup_sbox_0_output):(operation_274_5107_latch));
    assign operation_274_5106 = ((control_274_65)?(lookup_sbox_1_output):(operation_274_5106_latch));
    assign operation_274_5105 = ((control_274_65)?(lookup_sbox_2_output):(operation_274_5105_latch));
    assign operation_274_5104 = ((control_274_65)?(lookup_sbox_3_output):(operation_274_5104_latch));
    assign operation_274_5103 = ((control_274_65)?(lookup_sbox_4_output):(operation_274_5103_latch));
    assign operation_274_5102 = ((control_274_65)?(lookup_sbox_5_output):(operation_274_5102_latch));
    assign operation_274_5101 = ((control_274_65)?(lookup_sbox_6_output):(operation_274_5101_latch));
    assign operation_274_5100 = ((control_274_65)?(lookup_sbox_7_output):(operation_274_5100_latch));
    assign operation_274_5099 = ((control_274_65)?(lookup_sbox_8_output):(operation_274_5099_latch));
    assign operation_274_5098 = ((control_274_65)?(lookup_sbox_9_output):(operation_274_5098_latch));
    assign operation_274_5097 = ((control_274_65)?(lookup_sbox_10_output):(operation_274_5097_latch));
    assign operation_274_5096 = ((control_274_65)?(lookup_sbox_11_output):(operation_274_5096_latch));
    assign operation_274_5095 = ((control_274_65)?(lookup_sbox_12_output):(operation_274_5095_latch));
    assign operation_274_5094 = ((control_274_65)?(lookup_sbox_13_output):(operation_274_5094_latch));
    assign operation_274_5093 = ((control_274_65)?(lookup_sbox_14_output):(operation_274_5093_latch));
    assign operation_274_5092 = ((control_274_65)?(lookup_sbox_15_output):(operation_274_5092_latch));
    assign operation_274_1671 = ({(operation_274_1545[7:0])});
    assign operation_274_1535 = ({(operation_274_1505[7:0])});
    assign operation_274_1679 = ({(operation_274_1553[7:0])});
    assign operation_274_1655 = ({(operation_274_1529[7:0])});
    assign operation_274_4288 = (operation_274_4304);
    assign operation_274_4287 = (operation_274_4303);
    assign operation_274_4286 = (operation_274_4302);
    assign operation_274_4285 = (operation_274_4301);
    assign operation_274_4284 = (operation_274_4300);
    assign operation_274_4283 = (operation_274_4299);
    assign operation_274_4282 = (operation_274_4298);
    assign operation_274_4281 = (operation_274_4297);
    assign operation_274_4280 = (operation_274_4296);
    assign operation_274_4279 = (operation_274_4295);
    assign operation_274_4278 = (operation_274_4294);
    assign operation_274_4277 = (operation_274_4293);
    assign operation_274_4276 = (operation_274_4292);
    assign operation_274_4275 = (operation_274_4291);
    assign operation_274_4274 = (operation_274_4290);
    assign operation_274_4273 = (operation_274_4289);
    assign operation_274_1545 = (operation_274_1544);
    assign operation_274_1505 = (operation_274_1504);
    assign operation_274_1553 = (operation_274_1552);
    assign operation_274_1529 = (operation_274_1528);
    assign operation_274_4322 = ({(operation_274_4324[7:0])});
    assign operation_274_4321 = ({(operation_274_4325[7:0])});
    assign operation_274_4320 = ({(operation_274_4326[7:0])});
    assign operation_274_4319 = ({(operation_274_4327[7:0])});
    assign operation_274_4318 = ({(operation_274_4328[7:0])});
    assign operation_274_4317 = ({(operation_274_4329[7:0])});
    assign operation_274_4316 = ({(operation_274_4330[7:0])});
    assign operation_274_4315 = ({(operation_274_4331[7:0])});
    assign operation_274_4313 = ({(operation_274_4332[7:0])});
    assign operation_274_4312 = ({(operation_274_4333[7:0])});
    assign operation_274_4311 = ({(operation_274_4334[7:0])});
    assign operation_274_4310 = ({(operation_274_4335[7:0])});
    assign operation_274_4309 = ({(operation_274_4336[7:0])});
    assign operation_274_4308 = ({(operation_274_4337[7:0])});
    assign operation_274_4307 = ({(operation_274_4338[7:0])});
    assign operation_274_4305 = ({(operation_274_4339[7:0])});
    assign operation_274_1639 = ({(operation_274_1513[7:0])});
    assign operation_274_1503 = ({(operation_274_1473[7:0])});
    assign operation_274_1551 = ({(operation_274_1521[7:0])});
    assign operation_274_1623 = ({(operation_274_1497[7:0])});
    assign operation_274_4339 = (operation_274_4356);
    assign operation_274_4338 = (operation_274_4355);
    assign operation_274_4337 = (operation_274_4354);
    assign operation_274_4336 = (operation_274_4353);
    assign operation_274_4335 = (operation_274_4352);
    assign operation_274_4334 = (operation_274_4351);
    assign operation_274_4333 = (operation_274_4350);
    assign operation_274_4332 = (operation_274_4349);
    assign operation_274_4331 = (operation_274_4348);
    assign operation_274_4330 = (operation_274_4347);
    assign operation_274_4329 = (operation_274_4346);
    assign operation_274_4328 = (operation_274_4345);
    assign operation_274_4327 = (operation_274_4344);
    assign operation_274_4326 = (operation_274_4343);
    assign operation_274_4325 = (operation_274_4342);
    assign operation_274_4324 = (operation_274_4341);
    assign operation_274_1513 = (operation_274_1512);
    assign operation_274_1473 = (operation_274_1472);
    assign operation_274_1521 = (operation_274_1520);
    assign operation_274_1497 = (operation_274_1496);
    assign operation_274_4374 = ({(operation_274_4394[7:0])});
    assign operation_274_4373 = ({(operation_274_4393[7:0])});
    assign operation_274_4372 = ({(operation_274_4392[7:0])});
    assign operation_274_4371 = ({(operation_274_4391[7:0])});
    assign operation_274_4370 = ({(operation_274_4390[7:0])});
    assign operation_274_4369 = ({(operation_274_4389[7:0])});
    assign operation_274_4368 = ({(operation_274_4388[7:0])});
    assign operation_274_4367 = ({(operation_274_4387[7:0])});
    assign operation_274_4366 = ({(operation_274_4386[7:0])});
    assign operation_274_4365 = ({(operation_274_4385[7:0])});
    assign operation_274_4364 = ({(operation_274_4384[7:0])});
    assign operation_274_4363 = ({(operation_274_4383[7:0])});
    assign operation_274_4362 = ({(operation_274_4382[7:0])});
    assign operation_274_4361 = ({(operation_274_4381[7:0])});
    assign operation_274_4360 = ({(operation_274_4380[7:0])});
    assign operation_274_4359 = ({(operation_274_4379[7:0])});
    assign operation_274_1607 = ({(operation_274_1481[7:0])});
    assign operation_274_1471 = ({(operation_274_1441[7:0])});
    assign operation_274_1519 = ({(operation_274_1489[7:0])});
    assign operation_274_1591 = ({(operation_274_1465[7:0])});
    assign operation_274_4394 = (operation_274_4414);
    assign operation_274_4393 = (operation_274_4413);
    assign operation_274_4392 = (operation_274_4412);
    assign operation_274_4391 = (operation_274_4411);
    assign operation_274_4390 = (operation_274_4410);
    assign operation_274_4389 = (operation_274_4409);
    assign operation_274_4388 = (operation_274_4408);
    assign operation_274_4387 = (operation_274_4407);
    assign operation_274_4386 = (operation_274_4406);
    assign operation_274_4385 = (operation_274_4405);
    assign operation_274_4384 = (operation_274_4404);
    assign operation_274_4383 = (operation_274_4403);
    assign operation_274_4382 = (operation_274_4402);
    assign operation_274_4381 = (operation_274_4401);
    assign operation_274_4380 = (operation_274_4400);
    assign operation_274_4379 = (operation_274_4399);
    assign operation_274_1481 = (operation_274_1480);
    assign operation_274_1441 = (operation_274_1440);
    assign operation_274_1489 = (operation_274_1488);
    assign operation_274_1465 = (operation_274_1464);
    assign operation_274_4434 = ({(operation_274_4454[7:0])});
    assign operation_274_4433 = ({(operation_274_4453[7:0])});
    assign operation_274_4432 = ({(operation_274_4452[7:0])});
    assign operation_274_4431 = ({(operation_274_4451[7:0])});
    assign operation_274_4430 = ({(operation_274_4450[7:0])});
    assign operation_274_4429 = ({(operation_274_4449[7:0])});
    assign operation_274_4428 = ({(operation_274_4448[7:0])});
    assign operation_274_4427 = ({(operation_274_4447[7:0])});
    assign operation_274_4426 = ({(operation_274_4446[7:0])});
    assign operation_274_4425 = ({(operation_274_4445[7:0])});
    assign operation_274_4424 = ({(operation_274_4444[7:0])});
    assign operation_274_4423 = ({(operation_274_4443[7:0])});
    assign operation_274_4422 = ({(operation_274_4442[7:0])});
    assign operation_274_4421 = ({(operation_274_4441[7:0])});
    assign operation_274_4420 = ({(operation_274_4440[7:0])});
    assign operation_274_4419 = ({(operation_274_4439[7:0])});
    assign operation_274_1575 = ({(operation_274_1449[7:0])});
    assign operation_274_1439 = ({(operation_274_1433[7:0])});
    assign operation_274_1487 = ({(operation_274_1457[7:0])});
    assign operation_274_1463 = ({(operation_274_1423[7:0])});
    assign operation_274_4454 = (operation_274_4474);
    assign operation_274_4453 = (operation_274_4473);
    assign operation_274_4452 = (operation_274_4472);
    assign operation_274_4451 = (operation_274_4471);
    assign operation_274_4450 = (operation_274_4470);
    assign operation_274_4449 = (operation_274_4469);
    assign operation_274_4448 = (operation_274_4468);
    assign operation_274_4447 = (operation_274_4467);
    assign operation_274_4446 = (operation_274_4466);
    assign operation_274_4445 = (operation_274_4465);
    assign operation_274_4444 = (operation_274_4464);
    assign operation_274_4443 = (operation_274_4463);
    assign operation_274_4442 = (operation_274_4462);
    assign operation_274_4441 = (operation_274_4461);
    assign operation_274_4440 = (operation_274_4460);
    assign operation_274_4439 = (operation_274_4459);
    assign operation_274_5164 = ({(operation_274_5181[7:0])});
    assign operation_274_1449 = (operation_274_1448);
    assign operation_274_1433 = (operation_274_1432);
    assign operation_274_1457 = (operation_274_1456);
    assign operation_274_1423 = ((control_274_50)?(lookup_sbox_1_output):(operation_274_1423_latch));
    assign operation_274_5181 = (operation_274_5198);
    assign operation_274_1447 = ({(operation_274_1413[7:0])});
    assign operation_274_1428 = ({(operation_274_1408[7:0])});
    assign operation_274_1455 = ({(operation_274_1418[7:0])});
    assign operation_274_4502 = ({(operation_274_4557[7:0])});
    assign operation_274_4501 = ({(operation_274_4524[7:0])});
    assign operation_274_4500 = ({(operation_274_4558[7:0])});
    assign operation_274_4499 = ({(operation_274_4523[7:0])});
    assign operation_274_5234 = ({(operation_274_5254[7:0])});
    assign operation_274_5233 = ({(operation_274_5253[7:0])});
    assign operation_274_5216 = ({(operation_274_5236[7:0])});
    assign operation_274_5215 = ({(operation_274_5235[7:0])});
    assign operation_274_1418 = ((control_274_50)?(lookup_sbox_0_output):(operation_274_1418_latch));
    assign operation_274_1408 = ((control_274_49)?(lookup_sbox_0_output):(operation_274_1408_latch));
    assign operation_274_1413 = ((control_274_49)?(lookup_sbox_1_output):(operation_274_1413_latch));
    assign operation_274_4558 = (operation_274_4582);
    assign operation_274_4557 = (operation_274_4581);
    assign operation_274_4524 = (operation_274_4564);
    assign operation_274_4523 = (operation_274_4563);
    assign operation_274_5254 = (operation_274_5274);
    assign operation_274_5253 = (operation_274_5273);
    assign operation_274_5236 = (operation_274_5256);
    assign operation_274_5235 = (operation_274_5255);
    assign operation_274_4580 = ({(operation_274_4604[7:0])});
    assign operation_274_4579 = ({(operation_274_4603[7:0])});
    assign operation_274_4578 = ({(operation_274_4602[7:0])});
    assign operation_274_4577 = ({(operation_274_4601[7:0])});
    assign operation_274_4576 = ({(operation_274_4600[7:0])});
    assign operation_274_4575 = ({(operation_274_4599[7:0])});
    assign operation_274_4574 = ({(operation_274_4598[7:0])});
    assign operation_274_4573 = ({(operation_274_4597[7:0])});
    assign operation_274_4572 = ({(operation_274_4596[7:0])});
    assign operation_274_4571 = ({(operation_274_4595[7:0])});
    assign operation_274_4570 = ({(operation_274_4594[7:0])});
    assign operation_274_4569 = ({(operation_274_4593[7:0])});
    assign operation_274_4568 = ({(operation_274_4592[7:0])});
    assign operation_274_4567 = ({(operation_274_4591[7:0])});
    assign operation_274_4566 = ({(operation_274_4590[7:0])});
    assign operation_274_4565 = ({(operation_274_4589[7:0])});
    assign operation_274_4604 = (operation_274_4627);
    assign operation_274_4603 = (operation_274_4612);
    assign operation_274_4602 = (operation_274_4626);
    assign operation_274_4601 = (operation_274_4625);
    assign operation_274_4600 = (operation_274_4624);
    assign operation_274_4599 = (operation_274_4613);
    assign operation_274_4598 = (operation_274_4623);
    assign operation_274_4597 = (operation_274_4622);
    assign operation_274_4596 = (operation_274_4621);
    assign operation_274_4595 = (operation_274_4620);
    assign operation_274_4594 = (operation_274_4619);
    assign operation_274_4593 = (operation_274_4618);
    assign operation_274_4592 = (operation_274_4617);
    assign operation_274_4591 = (operation_274_4616);
    assign operation_274_4590 = (operation_274_4615);
    assign operation_274_4589 = (operation_274_4614);
    assign operation_274_5294 = ({(operation_274_5314[7:0])});
    assign operation_274_5293 = ({(operation_274_5313[7:0])});
    assign operation_274_5276 = ({(operation_274_5296[7:0])});
    assign operation_274_5275 = ({(operation_274_5295[7:0])});
    assign operation_274_5314 = (operation_274_5334);
    assign operation_274_5313 = (operation_274_5333);
    assign operation_274_5296 = (operation_274_5316);
    assign operation_274_5295 = (operation_274_5315);
    assign operation_274_4649 = ({(operation_274_4676[7:0])});
    assign operation_274_4648 = ({(operation_274_4671[7:0])});
    assign operation_274_4647 = ({(operation_274_4672[7:0])});
    assign operation_274_4646 = ({(operation_274_4675[7:0])});
    assign operation_274_4645 = ({(operation_274_4678[7:0])});
    assign operation_274_4644 = ({(operation_274_4673[7:0])});
    assign operation_274_4643 = ({(operation_274_4674[7:0])});
    assign operation_274_4642 = ({(operation_274_4677[7:0])});
    assign operation_274_4641 = ({(operation_274_4668[7:0])});
    assign operation_274_4640 = ({(operation_274_4663[7:0])});
    assign operation_274_4639 = ({(operation_274_4666[7:0])});
    assign operation_274_4638 = ({(operation_274_4669[7:0])});
    assign operation_274_4637 = ({(operation_274_4664[7:0])});
    assign operation_274_4636 = ({(operation_274_4667[7:0])});
    assign operation_274_4635 = ({(operation_274_4670[7:0])});
    assign operation_274_4634 = ({(operation_274_4665[7:0])});
    assign operation_274_4678 = ((control_274_56)?(lookup_sbox_0_output):(operation_274_4678_latch));
    assign operation_274_4677 = ((control_274_56)?(lookup_sbox_1_output):(operation_274_4677_latch));
    assign operation_274_4676 = ((control_274_56)?(lookup_sbox_2_output):(operation_274_4676_latch));
    assign operation_274_4675 = ((control_274_56)?(lookup_sbox_3_output):(operation_274_4675_latch));
    assign operation_274_4674 = ((control_274_56)?(lookup_sbox_4_output):(operation_274_4674_latch));
    assign operation_274_4673 = ((control_274_56)?(lookup_sbox_5_output):(operation_274_4673_latch));
    assign operation_274_4672 = ((control_274_56)?(lookup_sbox_6_output):(operation_274_4672_latch));
    assign operation_274_4671 = ((control_274_56)?(lookup_sbox_7_output):(operation_274_4671_latch));
    assign operation_274_4670 = ((control_274_56)?(lookup_sbox_8_output):(operation_274_4670_latch));
    assign operation_274_4669 = ((control_274_56)?(lookup_sbox_9_output):(operation_274_4669_latch));
    assign operation_274_4668 = ((control_274_56)?(lookup_sbox_10_output):(operation_274_4668_latch));
    assign operation_274_4667 = ((control_274_56)?(lookup_sbox_11_output):(operation_274_4667_latch));
    assign operation_274_4666 = ((control_274_56)?(lookup_sbox_12_output):(operation_274_4666_latch));
    assign operation_274_4665 = ((control_274_56)?(lookup_sbox_13_output):(operation_274_4665_latch));
    assign operation_274_4664 = ((control_274_56)?(lookup_sbox_14_output):(operation_274_4664_latch));
    assign operation_274_4663 = ((control_274_56)?(lookup_sbox_15_output):(operation_274_4663_latch));
    assign operation_274_5354 = ({(operation_274_5378[7:0])});
    assign operation_274_5353 = ({(operation_274_5377[7:0])});
    assign operation_274_5336 = ({(operation_274_5356[7:0])});
    assign operation_274_5335 = ({(operation_274_5355[7:0])});
    assign operation_274_3859 = (operation_274_3875);
    assign operation_274_3858 = (operation_274_3874);
    assign operation_274_3857 = (operation_274_3873);
    assign operation_274_3856 = (operation_274_3872);
    assign operation_274_3855 = (operation_274_3871);
    assign operation_274_3854 = (operation_274_3870);
    assign operation_274_3853 = (operation_274_3869);
    assign operation_274_3852 = (operation_274_3868);
    assign operation_274_3851 = (operation_274_3867);
    assign operation_274_3850 = (operation_274_3866);
    assign operation_274_3849 = (operation_274_3865);
    assign operation_274_3848 = (operation_274_3864);
    assign operation_274_3847 = (operation_274_3863);
    assign operation_274_3846 = (operation_274_3862);
    assign operation_274_3845 = (operation_274_3861);
    assign operation_274_3844 = (operation_274_3860);
    assign operation_274_5378 = (operation_274_5418);
    assign operation_274_5377 = (operation_274_5417);
    assign operation_274_5356 = (operation_274_5380);
    assign operation_274_5355 = (operation_274_5379);
    assign operation_274_3893 = ({(operation_274_3895[7:0])});
    assign operation_274_3892 = ({(operation_274_3896[7:0])});
    assign operation_274_3891 = ({(operation_274_3897[7:0])});
    assign operation_274_3890 = ({(operation_274_3898[7:0])});
    assign operation_274_3889 = ({(operation_274_3899[7:0])});
    assign operation_274_3888 = ({(operation_274_3900[7:0])});
    assign operation_274_3887 = ({(operation_274_3901[7:0])});
    assign operation_274_3886 = ({(operation_274_3902[7:0])});
    assign operation_274_3884 = ({(operation_274_3903[7:0])});
    assign operation_274_3883 = ({(operation_274_3904[7:0])});
    assign operation_274_3882 = ({(operation_274_3905[7:0])});
    assign operation_274_3881 = ({(operation_274_3906[7:0])});
    assign operation_274_3880 = ({(operation_274_3907[7:0])});
    assign operation_274_3879 = ({(operation_274_3908[7:0])});
    assign operation_274_3878 = ({(operation_274_3909[7:0])});
    assign operation_274_3876 = ({(operation_274_3910[7:0])});
    assign operation_274_5442 = ({(operation_274_5467[7:0])});
    assign operation_274_5441 = ({(operation_274_5466[7:0])});
    assign operation_274_5420 = ({(operation_274_5465[7:0])});
    assign operation_274_5419 = ({(operation_274_5444[7:0])});
    assign operation_274_3910 = (operation_274_3927);
    assign operation_274_3909 = (operation_274_3926);
    assign operation_274_3908 = (operation_274_3925);
    assign operation_274_3907 = (operation_274_3924);
    assign operation_274_3906 = (operation_274_3923);
    assign operation_274_3905 = (operation_274_3922);
    assign operation_274_3904 = (operation_274_3921);
    assign operation_274_3903 = (operation_274_3920);
    assign operation_274_3902 = (operation_274_3919);
    assign operation_274_3901 = (operation_274_3918);
    assign operation_274_3900 = (operation_274_3917);
    assign operation_274_3899 = (operation_274_3916);
    assign operation_274_3898 = (operation_274_3915);
    assign operation_274_3897 = (operation_274_3914);
    assign operation_274_3896 = (operation_274_3913);
    assign operation_274_3895 = (operation_274_3912);
    assign operation_274_5467 = (operation_274_5488);
    assign operation_274_5466 = (operation_274_5487);
    assign operation_274_5465 = (operation_274_5486);
    assign operation_274_5444 = (operation_274_5469);
    assign operation_274_3945 = ({(operation_274_3965[7:0])});
    assign operation_274_3944 = ({(operation_274_3964[7:0])});
    assign operation_274_3943 = ({(operation_274_3963[7:0])});
    assign operation_274_3942 = ({(operation_274_3962[7:0])});
    assign operation_274_3941 = ({(operation_274_3961[7:0])});
    assign operation_274_3940 = ({(operation_274_3960[7:0])});
    assign operation_274_3939 = ({(operation_274_3959[7:0])});
    assign operation_274_3938 = ({(operation_274_3958[7:0])});
    assign operation_274_3937 = ({(operation_274_3957[7:0])});
    assign operation_274_3936 = ({(operation_274_3956[7:0])});
    assign operation_274_3935 = ({(operation_274_3955[7:0])});
    assign operation_274_3934 = ({(operation_274_3954[7:0])});
    assign operation_274_3933 = ({(operation_274_3953[7:0])});
    assign operation_274_3932 = ({(operation_274_3952[7:0])});
    assign operation_274_3931 = ({(operation_274_3951[7:0])});
    assign operation_274_3930 = ({(operation_274_3950[7:0])});
    assign operation_274_5510 = ({(operation_274_5519[7:0])});
    assign operation_274_5509 = ({(operation_274_5520[7:0])});
    assign operation_274_5508 = ({(operation_274_5537[7:0])});
    assign operation_274_5491 = ({(operation_274_5538[7:0])});
    assign operation_274_3965 = (operation_274_3985);
    assign operation_274_3964 = (operation_274_3984);
    assign operation_274_3963 = (operation_274_3983);
    assign operation_274_3962 = (operation_274_3982);
    assign operation_274_3961 = (operation_274_3981);
    assign operation_274_3960 = (operation_274_3980);
    assign operation_274_3959 = (operation_274_3979);
    assign operation_274_3958 = (operation_274_3978);
    assign operation_274_3957 = (operation_274_3977);
    assign operation_274_3956 = (operation_274_3976);
    assign operation_274_3955 = (operation_274_3975);
    assign operation_274_3954 = (operation_274_3974);
    assign operation_274_3953 = (operation_274_3973);
    assign operation_274_3952 = (operation_274_3972);
    assign operation_274_3951 = (operation_274_3971);
    assign operation_274_3950 = (operation_274_3970);
    assign operation_274_4805 = ({(operation_274_4825[7:0])});
    assign operation_274_4804 = ({(operation_274_4824[7:0])});
    assign operation_274_4786 = ({(operation_274_4806[7:0])});
    assign operation_274_4735 = ({(operation_274_4752[7:0])});
    assign operation_274_5538 = ((control_274_44)?(lookup_sbox_2_output):(operation_274_5538_latch));
    assign operation_274_5537 = ((control_274_44)?(lookup_sbox_0_output):(operation_274_5537_latch));
    assign operation_274_5520 = ((control_274_44)?(lookup_sbox_1_output):(operation_274_5520_latch));
    assign operation_274_5519 = ((control_274_45)?(lookup_sbox_0_output):(operation_274_5519_latch));
    assign operation_274_4825 = (operation_274_4845);
    assign operation_274_4824 = (operation_274_4844);
    assign operation_274_4806 = (operation_274_4826);
    assign operation_274_4752 = (operation_274_4769);
    assign operation_274_4005 = ({(operation_274_4025[7:0])});
    assign operation_274_4004 = ({(operation_274_4024[7:0])});
    assign operation_274_4003 = ({(operation_274_4023[7:0])});
    assign operation_274_4002 = ({(operation_274_4022[7:0])});
    assign operation_274_4001 = ({(operation_274_4021[7:0])});
    assign operation_274_4000 = ({(operation_274_4020[7:0])});
    assign operation_274_3999 = ({(operation_274_4019[7:0])});
    assign operation_274_3998 = ({(operation_274_4018[7:0])});
    assign operation_274_3997 = ({(operation_274_4017[7:0])});
    assign operation_274_3996 = ({(operation_274_4016[7:0])});
    assign operation_274_3995 = ({(operation_274_4015[7:0])});
    assign operation_274_3994 = ({(operation_274_4014[7:0])});
    assign operation_274_3993 = ({(operation_274_4013[7:0])});
    assign operation_274_3992 = ({(operation_274_4012[7:0])});
    assign operation_274_3991 = ({(operation_274_4011[7:0])});
    assign operation_274_3990 = ({(operation_274_4010[7:0])});
    assign operation_274_4025 = (operation_274_4045);
    assign operation_274_4024 = (operation_274_4044);
    assign operation_274_4023 = (operation_274_4043);
    assign operation_274_4022 = (operation_274_4042);
    assign operation_274_4021 = (operation_274_4041);
    assign operation_274_4020 = (operation_274_4040);
    assign operation_274_4019 = (operation_274_4039);
    assign operation_274_4018 = (operation_274_4038);
    assign operation_274_4017 = (operation_274_4037);
    assign operation_274_4016 = (operation_274_4036);
    assign operation_274_4015 = (operation_274_4035);
    assign operation_274_4014 = (operation_274_4034);
    assign operation_274_4013 = (operation_274_4033);
    assign operation_274_4012 = (operation_274_4032);
    assign operation_274_4011 = (operation_274_4031);
    assign operation_274_4010 = (operation_274_4030);
    assign operation_274_4865 = ({(operation_274_4885[7:0])});
    assign operation_274_4864 = ({(operation_274_4884[7:0])});
    assign operation_274_4846 = ({(operation_274_4866[7:0])});
    assign operation_274_4787 = ({(operation_274_4807[7:0])});
    assign operation_274_4885 = (operation_274_4905);
    assign operation_274_4884 = (operation_274_4904);
    assign operation_274_4866 = (operation_274_4886);
    assign operation_274_4807 = (operation_274_4827);
    assign operation_274_4073 = ({(operation_274_4128[7:0])});
    assign operation_274_4072 = ({(operation_274_4095[7:0])});
    assign operation_274_4071 = ({(operation_274_4129[7:0])});
    assign operation_274_4070 = ({(operation_274_4094[7:0])});
    assign operation_274_4925 = ({(operation_274_4949[7:0])});
    assign operation_274_4924 = ({(operation_274_4948[7:0])});
    assign operation_274_4906 = ({(operation_274_4926[7:0])});
    assign operation_274_4847 = ({(operation_274_4867[7:0])});
    assign operation_274_4129 = (operation_274_4153);
    assign operation_274_4128 = (operation_274_4152);
    assign operation_274_4095 = (operation_274_4135);
    assign operation_274_4094 = (operation_274_4134);
    assign operation_274_4949 = (operation_274_4989);
    assign operation_274_4948 = (operation_274_4988);
    assign operation_274_4926 = (operation_274_4950);
    assign operation_274_4867 = (operation_274_4887);
    assign operation_274_4151 = ({(operation_274_4175[7:0])});
    assign operation_274_4150 = ({(operation_274_4174[7:0])});
    assign operation_274_4149 = ({(operation_274_4173[7:0])});
    assign operation_274_4148 = ({(operation_274_4172[7:0])});
    assign operation_274_4147 = ({(operation_274_4171[7:0])});
    assign operation_274_4146 = ({(operation_274_4170[7:0])});
    assign operation_274_4145 = ({(operation_274_4169[7:0])});
    assign operation_274_4144 = ({(operation_274_4168[7:0])});
    assign operation_274_4143 = ({(operation_274_4167[7:0])});
    assign operation_274_4142 = ({(operation_274_4166[7:0])});
    assign operation_274_4141 = ({(operation_274_4165[7:0])});
    assign operation_274_4140 = ({(operation_274_4164[7:0])});
    assign operation_274_4139 = ({(operation_274_4163[7:0])});
    assign operation_274_4138 = ({(operation_274_4162[7:0])});
    assign operation_274_4137 = ({(operation_274_4161[7:0])});
    assign operation_274_4136 = ({(operation_274_4160[7:0])});
    assign operation_274_4175 = (operation_274_4198);
    assign operation_274_4174 = (operation_274_4183);
    assign operation_274_4173 = (operation_274_4197);
    assign operation_274_4172 = (operation_274_4196);
    assign operation_274_4171 = (operation_274_4195);
    assign operation_274_4170 = (operation_274_4184);
    assign operation_274_4169 = (operation_274_4194);
    assign operation_274_4168 = (operation_274_4193);
    assign operation_274_4167 = (operation_274_4192);
    assign operation_274_4166 = (operation_274_4191);
    assign operation_274_4165 = (operation_274_4190);
    assign operation_274_4164 = (operation_274_4189);
    assign operation_274_4163 = (operation_274_4188);
    assign operation_274_4162 = (operation_274_4187);
    assign operation_274_4161 = (operation_274_4186);
    assign operation_274_4160 = (operation_274_4185);
    assign operation_274_5013 = ({(operation_274_5038[7:0])});
    assign operation_274_5012 = ({(operation_274_5037[7:0])});
    assign operation_274_4990 = ({(operation_274_5015[7:0])});
    assign operation_274_4907 = ({(operation_274_4927[7:0])});
    assign operation_274_5038 = (operation_274_5059);
    assign operation_274_5037 = (operation_274_5058);
    assign operation_274_5015 = (operation_274_5040);
    assign operation_274_4927 = (operation_274_4951);
    assign operation_274_4220 = ({(operation_274_4247[7:0])});
    assign operation_274_4219 = ({(operation_274_4242[7:0])});
    assign operation_274_4218 = ({(operation_274_4243[7:0])});
    assign operation_274_4217 = ({(operation_274_4246[7:0])});
    assign operation_274_4216 = ({(operation_274_4249[7:0])});
    assign operation_274_4215 = ({(operation_274_4244[7:0])});
    assign operation_274_4214 = ({(operation_274_4245[7:0])});
    assign operation_274_4213 = ({(operation_274_4248[7:0])});
    assign operation_274_4212 = ({(operation_274_4239[7:0])});
    assign operation_274_4211 = ({(operation_274_4234[7:0])});
    assign operation_274_4210 = ({(operation_274_4237[7:0])});
    assign operation_274_4209 = ({(operation_274_4240[7:0])});
    assign operation_274_4208 = ({(operation_274_4235[7:0])});
    assign operation_274_4207 = ({(operation_274_4238[7:0])});
    assign operation_274_4206 = ({(operation_274_4241[7:0])});
    assign operation_274_4205 = ({(operation_274_4236[7:0])});
    assign operation_274_4249 = ((control_274_47)?(lookup_sbox_0_output):(operation_274_4249_latch));
    assign operation_274_4248 = ((control_274_47)?(lookup_sbox_1_output):(operation_274_4248_latch));
    assign operation_274_4247 = ((control_274_47)?(lookup_sbox_2_output):(operation_274_4247_latch));
    assign operation_274_4246 = ((control_274_47)?(lookup_sbox_3_output):(operation_274_4246_latch));
    assign operation_274_4245 = ((control_274_47)?(lookup_sbox_4_output):(operation_274_4245_latch));
    assign operation_274_4244 = ((control_274_47)?(lookup_sbox_5_output):(operation_274_4244_latch));
    assign operation_274_4243 = ((control_274_47)?(lookup_sbox_6_output):(operation_274_4243_latch));
    assign operation_274_4242 = ((control_274_47)?(lookup_sbox_7_output):(operation_274_4242_latch));
    assign operation_274_4241 = ((control_274_47)?(lookup_sbox_8_output):(operation_274_4241_latch));
    assign operation_274_4240 = ((control_274_47)?(lookup_sbox_9_output):(operation_274_4240_latch));
    assign operation_274_4239 = ((control_274_47)?(lookup_sbox_10_output):(operation_274_4239_latch));
    assign operation_274_4238 = ((control_274_47)?(lookup_sbox_11_output):(operation_274_4238_latch));
    assign operation_274_4237 = ((control_274_47)?(lookup_sbox_12_output):(operation_274_4237_latch));
    assign operation_274_4236 = ((control_274_47)?(lookup_sbox_13_output):(operation_274_4236_latch));
    assign operation_274_4235 = ((control_274_47)?(lookup_sbox_14_output):(operation_274_4235_latch));
    assign operation_274_4234 = ((control_274_47)?(lookup_sbox_15_output):(operation_274_4234_latch));
    assign operation_274_5081 = ({(operation_274_5090[7:0])});
    assign operation_274_5080 = ({(operation_274_5091[7:0])});
    assign operation_274_5062 = ({(operation_274_5109[7:0])});
    assign operation_274_4991 = ({(operation_274_5036[7:0])});
    assign operation_274_3430 = (operation_274_3446);
    assign operation_274_3429 = (operation_274_3445);
    assign operation_274_3428 = (operation_274_3444);
    assign operation_274_3427 = (operation_274_3443);
    assign operation_274_3426 = (operation_274_3442);
    assign operation_274_3425 = (operation_274_3441);
    assign operation_274_3424 = (operation_274_3440);
    assign operation_274_3423 = (operation_274_3439);
    assign operation_274_3422 = (operation_274_3438);
    assign operation_274_3421 = (operation_274_3437);
    assign operation_274_3420 = (operation_274_3436);
    assign operation_274_3419 = (operation_274_3435);
    assign operation_274_3418 = (operation_274_3434);
    assign operation_274_3417 = (operation_274_3433);
    assign operation_274_3416 = (operation_274_3432);
    assign operation_274_3415 = (operation_274_3431);
    assign operation_274_4376 = ({(operation_274_4396[7:0])});
    assign operation_274_4357 = ({(operation_274_4377[7:0])});
    assign operation_274_4306 = ({(operation_274_4323[7:0])});
    assign operation_274_5109 = ((control_274_39)?(lookup_sbox_1_output):(operation_274_5109_latch));
    assign operation_274_5091 = ((control_274_39)?(lookup_sbox_2_output):(operation_274_5091_latch));
    assign operation_274_5090 = ((control_274_39)?(lookup_sbox_3_output):(operation_274_5090_latch));
    assign operation_274_5036 = (operation_274_5057);
    assign operation_274_4396 = (operation_274_4416);
    assign operation_274_4377 = (operation_274_4397);
    assign operation_274_4323 = (operation_274_4340);
    assign operation_274_3464 = ({(operation_274_3466[7:0])});
    assign operation_274_3463 = ({(operation_274_3467[7:0])});
    assign operation_274_3462 = ({(operation_274_3468[7:0])});
    assign operation_274_3461 = ({(operation_274_3469[7:0])});
    assign operation_274_3460 = ({(operation_274_3470[7:0])});
    assign operation_274_3459 = ({(operation_274_3471[7:0])});
    assign operation_274_3458 = ({(operation_274_3472[7:0])});
    assign operation_274_3457 = ({(operation_274_3473[7:0])});
    assign operation_274_3455 = ({(operation_274_3474[7:0])});
    assign operation_274_3454 = ({(operation_274_3475[7:0])});
    assign operation_274_3453 = ({(operation_274_3476[7:0])});
    assign operation_274_3452 = ({(operation_274_3477[7:0])});
    assign operation_274_3451 = ({(operation_274_3478[7:0])});
    assign operation_274_3450 = ({(operation_274_3479[7:0])});
    assign operation_274_3449 = ({(operation_274_3480[7:0])});
    assign operation_274_3447 = ({(operation_274_3481[7:0])});
    assign operation_274_5079 = ({(operation_274_5108[7:0])});
    assign operation_274_3481 = (operation_274_3498);
    assign operation_274_3480 = (operation_274_3497);
    assign operation_274_3479 = (operation_274_3496);
    assign operation_274_3478 = (operation_274_3495);
    assign operation_274_3477 = (operation_274_3494);
    assign operation_274_3476 = (operation_274_3493);
    assign operation_274_3475 = (operation_274_3492);
    assign operation_274_3474 = (operation_274_3491);
    assign operation_274_3473 = (operation_274_3490);
    assign operation_274_3472 = (operation_274_3489);
    assign operation_274_3471 = (operation_274_3488);
    assign operation_274_3470 = (operation_274_3487);
    assign operation_274_3469 = (operation_274_3486);
    assign operation_274_3468 = (operation_274_3485);
    assign operation_274_3467 = (operation_274_3484);
    assign operation_274_3466 = (operation_274_3483);
    assign operation_274_4436 = ({(operation_274_4456[7:0])});
    assign operation_274_4417 = ({(operation_274_4437[7:0])});
    assign operation_274_4375 = ({(operation_274_4395[7:0])});
    assign operation_274_4358 = ({(operation_274_4378[7:0])});
    assign operation_274_5108 = ((control_274_39)?(lookup_sbox_0_output):(operation_274_5108_latch));
    assign operation_274_4456 = (operation_274_4476);
    assign operation_274_4437 = (operation_274_4457);
    assign operation_274_4395 = (operation_274_4415);
    assign operation_274_4378 = (operation_274_4398);
    assign operation_274_3516 = ({(operation_274_3536[7:0])});
    assign operation_274_3515 = ({(operation_274_3535[7:0])});
    assign operation_274_3514 = ({(operation_274_3534[7:0])});
    assign operation_274_3513 = ({(operation_274_3533[7:0])});
    assign operation_274_3512 = ({(operation_274_3532[7:0])});
    assign operation_274_3511 = ({(operation_274_3531[7:0])});
    assign operation_274_3510 = ({(operation_274_3530[7:0])});
    assign operation_274_3509 = ({(operation_274_3529[7:0])});
    assign operation_274_3508 = ({(operation_274_3528[7:0])});
    assign operation_274_3507 = ({(operation_274_3527[7:0])});
    assign operation_274_3506 = ({(operation_274_3526[7:0])});
    assign operation_274_3505 = ({(operation_274_3525[7:0])});
    assign operation_274_3504 = ({(operation_274_3524[7:0])});
    assign operation_274_3503 = ({(operation_274_3523[7:0])});
    assign operation_274_3502 = ({(operation_274_3522[7:0])});
    assign operation_274_3501 = ({(operation_274_3521[7:0])});
    assign operation_274_3536 = (operation_274_3556);
    assign operation_274_3535 = (operation_274_3555);
    assign operation_274_3534 = (operation_274_3554);
    assign operation_274_3533 = (operation_274_3553);
    assign operation_274_3532 = (operation_274_3552);
    assign operation_274_3531 = (operation_274_3551);
    assign operation_274_3530 = (operation_274_3550);
    assign operation_274_3529 = (operation_274_3549);
    assign operation_274_3528 = (operation_274_3548);
    assign operation_274_3527 = (operation_274_3547);
    assign operation_274_3526 = (operation_274_3546);
    assign operation_274_3525 = (operation_274_3545);
    assign operation_274_3524 = (operation_274_3544);
    assign operation_274_3523 = (operation_274_3543);
    assign operation_274_3522 = (operation_274_3542);
    assign operation_274_3521 = (operation_274_3541);
    assign operation_274_4496 = ({(operation_274_4520[7:0])});
    assign operation_274_4477 = ({(operation_274_4497[7:0])});
    assign operation_274_4435 = ({(operation_274_4455[7:0])});
    assign operation_274_4418 = ({(operation_274_4438[7:0])});
    assign operation_274_4520 = (operation_274_4560);
    assign operation_274_4497 = (operation_274_4521);
    assign operation_274_4455 = (operation_274_4475);
    assign operation_274_4438 = (operation_274_4458);
    assign operation_274_3576 = ({(operation_274_3596[7:0])});
    assign operation_274_3575 = ({(operation_274_3595[7:0])});
    assign operation_274_3574 = ({(operation_274_3594[7:0])});
    assign operation_274_3573 = ({(operation_274_3593[7:0])});
    assign operation_274_3572 = ({(operation_274_3592[7:0])});
    assign operation_274_3571 = ({(operation_274_3591[7:0])});
    assign operation_274_3570 = ({(operation_274_3590[7:0])});
    assign operation_274_3569 = ({(operation_274_3589[7:0])});
    assign operation_274_3568 = ({(operation_274_3588[7:0])});
    assign operation_274_3567 = ({(operation_274_3587[7:0])});
    assign operation_274_3566 = ({(operation_274_3586[7:0])});
    assign operation_274_3565 = ({(operation_274_3585[7:0])});
    assign operation_274_3564 = ({(operation_274_3584[7:0])});
    assign operation_274_3563 = ({(operation_274_3583[7:0])});
    assign operation_274_3562 = ({(operation_274_3582[7:0])});
    assign operation_274_3561 = ({(operation_274_3581[7:0])});
    assign operation_274_3596 = (operation_274_3616);
    assign operation_274_3595 = (operation_274_3615);
    assign operation_274_3594 = (operation_274_3614);
    assign operation_274_3593 = (operation_274_3613);
    assign operation_274_3592 = (operation_274_3612);
    assign operation_274_3591 = (operation_274_3611);
    assign operation_274_3590 = (operation_274_3610);
    assign operation_274_3589 = (operation_274_3609);
    assign operation_274_3588 = (operation_274_3608);
    assign operation_274_3587 = (operation_274_3607);
    assign operation_274_3586 = (operation_274_3606);
    assign operation_274_3585 = (operation_274_3605);
    assign operation_274_3584 = (operation_274_3604);
    assign operation_274_3583 = (operation_274_3603);
    assign operation_274_3582 = (operation_274_3602);
    assign operation_274_3581 = (operation_274_3601);
    assign operation_274_4584 = ({(operation_274_4609[7:0])});
    assign operation_274_4561 = ({(operation_274_4586[7:0])});
    assign operation_274_4495 = ({(operation_274_4519[7:0])});
    assign operation_274_4478 = ({(operation_274_4498[7:0])});
    assign operation_274_4609 = (operation_274_4630);
    assign operation_274_4586 = (operation_274_4611);
    assign operation_274_4519 = (operation_274_4559);
    assign operation_274_4498 = (operation_274_4522);
    assign operation_274_3644 = ({(operation_274_3699[7:0])});
    assign operation_274_3643 = ({(operation_274_3666[7:0])});
    assign operation_274_3642 = ({(operation_274_3700[7:0])});
    assign operation_274_3641 = ({(operation_274_3665[7:0])});
    assign operation_274_4652 = ({(operation_274_4661[7:0])});
    assign operation_274_4633 = ({(operation_274_4680[7:0])});
    assign operation_274_4583 = ({(operation_274_4608[7:0])});
    assign operation_274_4562 = ({(operation_274_4607[7:0])});
    assign operation_274_3700 = (operation_274_3724);
    assign operation_274_3699 = (operation_274_3723);
    assign operation_274_3666 = (operation_274_3706);
    assign operation_274_3665 = (operation_274_3705);
    assign operation_274_3947 = ({(operation_274_3967[7:0])});
    assign operation_274_3877 = ({(operation_274_3894[7:0])});
    assign operation_274_4680 = ((control_274_33)?(lookup_sbox_2_output):(operation_274_4680_latch));
    assign operation_274_4661 = ((control_274_33)?(lookup_sbox_3_output):(operation_274_4661_latch));
    assign operation_274_4608 = (operation_274_4629);
    assign operation_274_4607 = (operation_274_4628);
    assign operation_274_3722 = ({(operation_274_3746[7:0])});
    assign operation_274_3721 = ({(operation_274_3745[7:0])});
    assign operation_274_3720 = ({(operation_274_3744[7:0])});
    assign operation_274_3719 = ({(operation_274_3743[7:0])});
    assign operation_274_3718 = ({(operation_274_3742[7:0])});
    assign operation_274_3717 = ({(operation_274_3741[7:0])});
    assign operation_274_3716 = ({(operation_274_3740[7:0])});
    assign operation_274_3715 = ({(operation_274_3739[7:0])});
    assign operation_274_3714 = ({(operation_274_3738[7:0])});
    assign operation_274_3713 = ({(operation_274_3737[7:0])});
    assign operation_274_3712 = ({(operation_274_3736[7:0])});
    assign operation_274_3711 = ({(operation_274_3735[7:0])});
    assign operation_274_3710 = ({(operation_274_3734[7:0])});
    assign operation_274_3709 = ({(operation_274_3733[7:0])});
    assign operation_274_3708 = ({(operation_274_3732[7:0])});
    assign operation_274_3707 = ({(operation_274_3731[7:0])});
    assign operation_274_3967 = (operation_274_3987);
    assign operation_274_3894 = (operation_274_3911);
    assign operation_274_3746 = (operation_274_3769);
    assign operation_274_3745 = (operation_274_3754);
    assign operation_274_3744 = (operation_274_3768);
    assign operation_274_3743 = (operation_274_3767);
    assign operation_274_3742 = (operation_274_3766);
    assign operation_274_3741 = (operation_274_3755);
    assign operation_274_3740 = (operation_274_3765);
    assign operation_274_3739 = (operation_274_3764);
    assign operation_274_3738 = (operation_274_3763);
    assign operation_274_3737 = (operation_274_3762);
    assign operation_274_3736 = (operation_274_3761);
    assign operation_274_3735 = (operation_274_3760);
    assign operation_274_3734 = (operation_274_3759);
    assign operation_274_3733 = (operation_274_3758);
    assign operation_274_3732 = (operation_274_3757);
    assign operation_274_3731 = (operation_274_3756);
    assign operation_274_4651 = ({(operation_274_4662[7:0])});
    assign operation_274_4650 = ({(operation_274_4679[7:0])});
    assign operation_274_4007 = ({(operation_274_4027[7:0])});
    assign operation_274_3946 = ({(operation_274_3966[7:0])});
    assign operation_274_3929 = ({(operation_274_3949[7:0])});
    assign operation_274_3928 = ({(operation_274_3948[7:0])});
    assign operation_274_4679 = ((control_274_33)?(lookup_sbox_0_output):(operation_274_4679_latch));
    assign operation_274_4662 = ((control_274_33)?(lookup_sbox_1_output):(operation_274_4662_latch));
    assign operation_274_3791 = ({(operation_274_3818[7:0])});
    assign operation_274_3790 = ({(operation_274_3813[7:0])});
    assign operation_274_3789 = ({(operation_274_3814[7:0])});
    assign operation_274_3788 = ({(operation_274_3817[7:0])});
    assign operation_274_3787 = ({(operation_274_3820[7:0])});
    assign operation_274_3786 = ({(operation_274_3815[7:0])});
    assign operation_274_3785 = ({(operation_274_3816[7:0])});
    assign operation_274_3784 = ({(operation_274_3819[7:0])});
    assign operation_274_3783 = ({(operation_274_3810[7:0])});
    assign operation_274_3782 = ({(operation_274_3805[7:0])});
    assign operation_274_3781 = ({(operation_274_3808[7:0])});
    assign operation_274_3780 = ({(operation_274_3811[7:0])});
    assign operation_274_3779 = ({(operation_274_3806[7:0])});
    assign operation_274_3778 = ({(operation_274_3809[7:0])});
    assign operation_274_3777 = ({(operation_274_3812[7:0])});
    assign operation_274_3776 = ({(operation_274_3807[7:0])});
    assign operation_274_4027 = (operation_274_4047);
    assign operation_274_3966 = (operation_274_3986);
    assign operation_274_3949 = (operation_274_3969);
    assign operation_274_3948 = (operation_274_3968);
    assign operation_274_3820 = ((control_274_38)?(lookup_sbox_0_output):(operation_274_3820_latch));
    assign operation_274_3819 = ((control_274_38)?(lookup_sbox_1_output):(operation_274_3819_latch));
    assign operation_274_3818 = ((control_274_38)?(lookup_sbox_2_output):(operation_274_3818_latch));
    assign operation_274_3817 = ((control_274_38)?(lookup_sbox_3_output):(operation_274_3817_latch));
    assign operation_274_3816 = ((control_274_38)?(lookup_sbox_4_output):(operation_274_3816_latch));
    assign operation_274_3815 = ((control_274_38)?(lookup_sbox_5_output):(operation_274_3815_latch));
    assign operation_274_3814 = ((control_274_38)?(lookup_sbox_6_output):(operation_274_3814_latch));
    assign operation_274_3813 = ((control_274_38)?(lookup_sbox_7_output):(operation_274_3813_latch));
    assign operation_274_3812 = ((control_274_38)?(lookup_sbox_8_output):(operation_274_3812_latch));
    assign operation_274_3811 = ((control_274_38)?(lookup_sbox_9_output):(operation_274_3811_latch));
    assign operation_274_3810 = ((control_274_38)?(lookup_sbox_10_output):(operation_274_3810_latch));
    assign operation_274_3809 = ((control_274_38)?(lookup_sbox_11_output):(operation_274_3809_latch));
    assign operation_274_3808 = ((control_274_38)?(lookup_sbox_12_output):(operation_274_3808_latch));
    assign operation_274_3807 = ((control_274_38)?(lookup_sbox_13_output):(operation_274_3807_latch));
    assign operation_274_3806 = ((control_274_38)?(lookup_sbox_14_output):(operation_274_3806_latch));
    assign operation_274_3805 = ((control_274_38)?(lookup_sbox_15_output):(operation_274_3805_latch));
    assign operation_274_3001 = (operation_274_3017);
    assign operation_274_3000 = (operation_274_3016);
    assign operation_274_2999 = (operation_274_3015);
    assign operation_274_2998 = (operation_274_3014);
    assign operation_274_2997 = (operation_274_3013);
    assign operation_274_2996 = (operation_274_3012);
    assign operation_274_2995 = (operation_274_3011);
    assign operation_274_2994 = (operation_274_3010);
    assign operation_274_2993 = (operation_274_3009);
    assign operation_274_2992 = (operation_274_3008);
    assign operation_274_2991 = (operation_274_3007);
    assign operation_274_2990 = (operation_274_3006);
    assign operation_274_2989 = (operation_274_3005);
    assign operation_274_2988 = (operation_274_3004);
    assign operation_274_2987 = (operation_274_3003);
    assign operation_274_2986 = (operation_274_3002);
    assign operation_274_4067 = ({(operation_274_4091[7:0])});
    assign operation_274_4006 = ({(operation_274_4026[7:0])});
    assign operation_274_3989 = ({(operation_274_4009[7:0])});
    assign operation_274_3988 = ({(operation_274_4008[7:0])});
    assign operation_274_4091 = (operation_274_4131);
    assign operation_274_4026 = (operation_274_4046);
    assign operation_274_4009 = (operation_274_4029);
    assign operation_274_4008 = (operation_274_4028);
    assign operation_274_3035 = ({(operation_274_3037[7:0])});
    assign operation_274_3034 = ({(operation_274_3038[7:0])});
    assign operation_274_3033 = ({(operation_274_3039[7:0])});
    assign operation_274_3032 = ({(operation_274_3040[7:0])});
    assign operation_274_3031 = ({(operation_274_3041[7:0])});
    assign operation_274_3030 = ({(operation_274_3042[7:0])});
    assign operation_274_3029 = ({(operation_274_3043[7:0])});
    assign operation_274_3028 = ({(operation_274_3044[7:0])});
    assign operation_274_3026 = ({(operation_274_3045[7:0])});
    assign operation_274_3025 = ({(operation_274_3046[7:0])});
    assign operation_274_3024 = ({(operation_274_3047[7:0])});
    assign operation_274_3023 = ({(operation_274_3048[7:0])});
    assign operation_274_3022 = ({(operation_274_3049[7:0])});
    assign operation_274_3021 = ({(operation_274_3050[7:0])});
    assign operation_274_3020 = ({(operation_274_3051[7:0])});
    assign operation_274_3018 = ({(operation_274_3052[7:0])});
    assign operation_274_3052 = (operation_274_3069);
    assign operation_274_3051 = (operation_274_3068);
    assign operation_274_3050 = (operation_274_3067);
    assign operation_274_3049 = (operation_274_3066);
    assign operation_274_3048 = (operation_274_3065);
    assign operation_274_3047 = (operation_274_3064);
    assign operation_274_3046 = (operation_274_3063);
    assign operation_274_3045 = (operation_274_3062);
    assign operation_274_3044 = (operation_274_3061);
    assign operation_274_3043 = (operation_274_3060);
    assign operation_274_3042 = (operation_274_3059);
    assign operation_274_3041 = (operation_274_3058);
    assign operation_274_3040 = (operation_274_3057);
    assign operation_274_3039 = (operation_274_3056);
    assign operation_274_3038 = (operation_274_3055);
    assign operation_274_3037 = (operation_274_3054);
    assign operation_274_4155 = ({(operation_274_4180[7:0])});
    assign operation_274_4066 = ({(operation_274_4090[7:0])});
    assign operation_274_4049 = ({(operation_274_4069[7:0])});
    assign operation_274_4048 = ({(operation_274_4068[7:0])});
    assign operation_274_4180 = (operation_274_4201);
    assign operation_274_4090 = (operation_274_4130);
    assign operation_274_4069 = (operation_274_4093);
    assign operation_274_4068 = (operation_274_4092);
    assign operation_274_3087 = ({(operation_274_3107[7:0])});
    assign operation_274_3086 = ({(operation_274_3106[7:0])});
    assign operation_274_3085 = ({(operation_274_3105[7:0])});
    assign operation_274_3084 = ({(operation_274_3104[7:0])});
    assign operation_274_3083 = ({(operation_274_3103[7:0])});
    assign operation_274_3082 = ({(operation_274_3102[7:0])});
    assign operation_274_3081 = ({(operation_274_3101[7:0])});
    assign operation_274_3080 = ({(operation_274_3100[7:0])});
    assign operation_274_3079 = ({(operation_274_3099[7:0])});
    assign operation_274_3078 = ({(operation_274_3098[7:0])});
    assign operation_274_3077 = ({(operation_274_3097[7:0])});
    assign operation_274_3076 = ({(operation_274_3096[7:0])});
    assign operation_274_3075 = ({(operation_274_3095[7:0])});
    assign operation_274_3074 = ({(operation_274_3094[7:0])});
    assign operation_274_3073 = ({(operation_274_3093[7:0])});
    assign operation_274_3072 = ({(operation_274_3092[7:0])});
    assign operation_274_3107 = (operation_274_3127);
    assign operation_274_3106 = (operation_274_3126);
    assign operation_274_3105 = (operation_274_3125);
    assign operation_274_3104 = (operation_274_3124);
    assign operation_274_3103 = (operation_274_3123);
    assign operation_274_3102 = (operation_274_3122);
    assign operation_274_3101 = (operation_274_3121);
    assign operation_274_3100 = (operation_274_3120);
    assign operation_274_3099 = (operation_274_3119);
    assign operation_274_3098 = (operation_274_3118);
    assign operation_274_3097 = (operation_274_3117);
    assign operation_274_3096 = (operation_274_3116);
    assign operation_274_3095 = (operation_274_3115);
    assign operation_274_3094 = (operation_274_3114);
    assign operation_274_3093 = (operation_274_3113);
    assign operation_274_3092 = (operation_274_3112);
    assign operation_274_4223 = ({(operation_274_4232[7:0])});
    assign operation_274_4154 = ({(operation_274_4179[7:0])});
    assign operation_274_4133 = ({(operation_274_4178[7:0])});
    assign operation_274_4132 = ({(operation_274_4157[7:0])});
    assign operation_274_3448 = ({(operation_274_3465[7:0])});
    assign operation_274_4232 = ((control_274_28)?(lookup_sbox_2_output):(operation_274_4232_latch));
    assign operation_274_4179 = (operation_274_4200);
    assign operation_274_4178 = (operation_274_4199);
    assign operation_274_4157 = (operation_274_4182);
    assign operation_274_3147 = ({(operation_274_3167[7:0])});
    assign operation_274_3146 = ({(operation_274_3166[7:0])});
    assign operation_274_3145 = ({(operation_274_3165[7:0])});
    assign operation_274_3144 = ({(operation_274_3164[7:0])});
    assign operation_274_3143 = ({(operation_274_3163[7:0])});
    assign operation_274_3142 = ({(operation_274_3162[7:0])});
    assign operation_274_3141 = ({(operation_274_3161[7:0])});
    assign operation_274_3140 = ({(operation_274_3160[7:0])});
    assign operation_274_3139 = ({(operation_274_3159[7:0])});
    assign operation_274_3138 = ({(operation_274_3158[7:0])});
    assign operation_274_3137 = ({(operation_274_3157[7:0])});
    assign operation_274_3136 = ({(operation_274_3156[7:0])});
    assign operation_274_3135 = ({(operation_274_3155[7:0])});
    assign operation_274_3134 = ({(operation_274_3154[7:0])});
    assign operation_274_3133 = ({(operation_274_3153[7:0])});
    assign operation_274_3132 = ({(operation_274_3152[7:0])});
    assign operation_274_3465 = (operation_274_3482);
    assign operation_274_3167 = (operation_274_3187);
    assign operation_274_3166 = (operation_274_3186);
    assign operation_274_3165 = (operation_274_3185);
    assign operation_274_3164 = (operation_274_3184);
    assign operation_274_3163 = (operation_274_3183);
    assign operation_274_3162 = (operation_274_3182);
    assign operation_274_3161 = (operation_274_3181);
    assign operation_274_3160 = (operation_274_3180);
    assign operation_274_3159 = (operation_274_3179);
    assign operation_274_3158 = (operation_274_3178);
    assign operation_274_3157 = (operation_274_3177);
    assign operation_274_3156 = (operation_274_3176);
    assign operation_274_3155 = (operation_274_3175);
    assign operation_274_3154 = (operation_274_3174);
    assign operation_274_3153 = (operation_274_3173);
    assign operation_274_3152 = (operation_274_3172);
    assign operation_274_4222 = ({(operation_274_4233[7:0])});
    assign operation_274_4221 = ({(operation_274_4250[7:0])});
    assign operation_274_4204 = ({(operation_274_4251[7:0])});
    assign operation_274_3518 = ({(operation_274_3538[7:0])});
    assign operation_274_3517 = ({(operation_274_3537[7:0])});
    assign operation_274_3500 = ({(operation_274_3520[7:0])});
    assign operation_274_3499 = ({(operation_274_3519[7:0])});
    assign operation_274_4251 = ((control_274_28)?(lookup_sbox_0_output):(operation_274_4251_latch));
    assign operation_274_4250 = ((control_274_27)?(lookup_sbox_0_output):(operation_274_4250_latch));
    assign operation_274_4233 = ((control_274_28)?(lookup_sbox_1_output):(operation_274_4233_latch));
    assign operation_274_3538 = (operation_274_3558);
    assign operation_274_3537 = (operation_274_3557);
    assign operation_274_3520 = (operation_274_3540);
    assign operation_274_3519 = (operation_274_3539);
    assign operation_274_3215 = ({(operation_274_3270[7:0])});
    assign operation_274_3214 = ({(operation_274_3237[7:0])});
    assign operation_274_3213 = ({(operation_274_3271[7:0])});
    assign operation_274_3212 = ({(operation_274_3236[7:0])});
    assign operation_274_3271 = (operation_274_3295);
    assign operation_274_3270 = (operation_274_3294);
    assign operation_274_3237 = (operation_274_3277);
    assign operation_274_3236 = (operation_274_3276);
    assign operation_274_3578 = ({(operation_274_3598[7:0])});
    assign operation_274_3577 = ({(operation_274_3597[7:0])});
    assign operation_274_3560 = ({(operation_274_3580[7:0])});
    assign operation_274_3559 = ({(operation_274_3579[7:0])});
    assign operation_274_3293 = ({(operation_274_3317[7:0])});
    assign operation_274_3292 = ({(operation_274_3316[7:0])});
    assign operation_274_3291 = ({(operation_274_3315[7:0])});
    assign operation_274_3290 = ({(operation_274_3314[7:0])});
    assign operation_274_3289 = ({(operation_274_3313[7:0])});
    assign operation_274_3288 = ({(operation_274_3312[7:0])});
    assign operation_274_3287 = ({(operation_274_3311[7:0])});
    assign operation_274_3286 = ({(operation_274_3310[7:0])});
    assign operation_274_3285 = ({(operation_274_3309[7:0])});
    assign operation_274_3284 = ({(operation_274_3308[7:0])});
    assign operation_274_3283 = ({(operation_274_3307[7:0])});
    assign operation_274_3282 = ({(operation_274_3306[7:0])});
    assign operation_274_3281 = ({(operation_274_3305[7:0])});
    assign operation_274_3280 = ({(operation_274_3304[7:0])});
    assign operation_274_3279 = ({(operation_274_3303[7:0])});
    assign operation_274_3278 = ({(operation_274_3302[7:0])});
    assign operation_274_3598 = (operation_274_3618);
    assign operation_274_3597 = (operation_274_3617);
    assign operation_274_3580 = (operation_274_3600);
    assign operation_274_3579 = (operation_274_3599);
    assign operation_274_3317 = (operation_274_3340);
    assign operation_274_3316 = (operation_274_3325);
    assign operation_274_3315 = (operation_274_3339);
    assign operation_274_3314 = (operation_274_3338);
    assign operation_274_3313 = (operation_274_3337);
    assign operation_274_3312 = (operation_274_3326);
    assign operation_274_3311 = (operation_274_3336);
    assign operation_274_3310 = (operation_274_3335);
    assign operation_274_3309 = (operation_274_3334);
    assign operation_274_3308 = (operation_274_3333);
    assign operation_274_3307 = (operation_274_3332);
    assign operation_274_3306 = (operation_274_3331);
    assign operation_274_3305 = (operation_274_3330);
    assign operation_274_3304 = (operation_274_3329);
    assign operation_274_3303 = (operation_274_3328);
    assign operation_274_3302 = (operation_274_3327);
    assign operation_274_3638 = ({(operation_274_3662[7:0])});
    assign operation_274_3637 = ({(operation_274_3661[7:0])});
    assign operation_274_3620 = ({(operation_274_3640[7:0])});
    assign operation_274_3619 = ({(operation_274_3639[7:0])});
    assign operation_274_3362 = ({(operation_274_3389[7:0])});
    assign operation_274_3361 = ({(operation_274_3384[7:0])});
    assign operation_274_3360 = ({(operation_274_3385[7:0])});
    assign operation_274_3359 = ({(operation_274_3388[7:0])});
    assign operation_274_3358 = ({(operation_274_3391[7:0])});
    assign operation_274_3357 = ({(operation_274_3386[7:0])});
    assign operation_274_3356 = ({(operation_274_3387[7:0])});
    assign operation_274_3355 = ({(operation_274_3390[7:0])});
    assign operation_274_3354 = ({(operation_274_3381[7:0])});
    assign operation_274_3353 = ({(operation_274_3376[7:0])});
    assign operation_274_3352 = ({(operation_274_3379[7:0])});
    assign operation_274_3351 = ({(operation_274_3382[7:0])});
    assign operation_274_3350 = ({(operation_274_3377[7:0])});
    assign operation_274_3349 = ({(operation_274_3380[7:0])});
    assign operation_274_3348 = ({(operation_274_3383[7:0])});
    assign operation_274_3347 = ({(operation_274_3378[7:0])});
    assign operation_274_3662 = (operation_274_3702);
    assign operation_274_3661 = (operation_274_3701);
    assign operation_274_3640 = (operation_274_3664);
    assign operation_274_3639 = (operation_274_3663);
    assign operation_274_3391 = ((control_274_29)?(lookup_sbox_0_output):(operation_274_3391_latch));
    assign operation_274_3390 = ((control_274_29)?(lookup_sbox_1_output):(operation_274_3390_latch));
    assign operation_274_3389 = ((control_274_29)?(lookup_sbox_2_output):(operation_274_3389_latch));
    assign operation_274_3388 = ((control_274_29)?(lookup_sbox_3_output):(operation_274_3388_latch));
    assign operation_274_3387 = ((control_274_29)?(lookup_sbox_4_output):(operation_274_3387_latch));
    assign operation_274_3386 = ((control_274_29)?(lookup_sbox_5_output):(operation_274_3386_latch));
    assign operation_274_3385 = ((control_274_29)?(lookup_sbox_6_output):(operation_274_3385_latch));
    assign operation_274_3384 = ((control_274_29)?(lookup_sbox_7_output):(operation_274_3384_latch));
    assign operation_274_3383 = ((control_274_29)?(lookup_sbox_8_output):(operation_274_3383_latch));
    assign operation_274_3382 = ((control_274_29)?(lookup_sbox_9_output):(operation_274_3382_latch));
    assign operation_274_3381 = ((control_274_29)?(lookup_sbox_10_output):(operation_274_3381_latch));
    assign operation_274_3380 = ((control_274_29)?(lookup_sbox_11_output):(operation_274_3380_latch));
    assign operation_274_3379 = ((control_274_29)?(lookup_sbox_12_output):(operation_274_3379_latch));
    assign operation_274_3378 = ((control_274_29)?(lookup_sbox_13_output):(operation_274_3378_latch));
    assign operation_274_3377 = ((control_274_29)?(lookup_sbox_14_output):(operation_274_3377_latch));
    assign operation_274_3376 = ((control_274_29)?(lookup_sbox_15_output):(operation_274_3376_latch));
    assign operation_274_2572 = (operation_274_2588);
    assign operation_274_2571 = (operation_274_2587);
    assign operation_274_2570 = (operation_274_2586);
    assign operation_274_2569 = (operation_274_2585);
    assign operation_274_2568 = (operation_274_2584);
    assign operation_274_2567 = (operation_274_2583);
    assign operation_274_2566 = (operation_274_2582);
    assign operation_274_2565 = (operation_274_2581);
    assign operation_274_2564 = (operation_274_2580);
    assign operation_274_2563 = (operation_274_2579);
    assign operation_274_2562 = (operation_274_2578);
    assign operation_274_2561 = (operation_274_2577);
    assign operation_274_2560 = (operation_274_2576);
    assign operation_274_2559 = (operation_274_2575);
    assign operation_274_2558 = (operation_274_2574);
    assign operation_274_2557 = (operation_274_2573);
    assign operation_274_3726 = ({(operation_274_3751[7:0])});
    assign operation_274_3725 = ({(operation_274_3750[7:0])});
    assign operation_274_3704 = ({(operation_274_3749[7:0])});
    assign operation_274_3703 = ({(operation_274_3728[7:0])});
    assign operation_274_3751 = (operation_274_3772);
    assign operation_274_3750 = (operation_274_3771);
    assign operation_274_3749 = (operation_274_3770);
    assign operation_274_3728 = (operation_274_3753);
    assign operation_274_2606 = ({(operation_274_2608[7:0])});
    assign operation_274_2605 = ({(operation_274_2609[7:0])});
    assign operation_274_2604 = ({(operation_274_2610[7:0])});
    assign operation_274_2603 = ({(operation_274_2611[7:0])});
    assign operation_274_2602 = ({(operation_274_2612[7:0])});
    assign operation_274_2601 = ({(operation_274_2613[7:0])});
    assign operation_274_2600 = ({(operation_274_2614[7:0])});
    assign operation_274_2599 = ({(operation_274_2615[7:0])});
    assign operation_274_2597 = ({(operation_274_2616[7:0])});
    assign operation_274_2596 = ({(operation_274_2617[7:0])});
    assign operation_274_2595 = ({(operation_274_2618[7:0])});
    assign operation_274_2594 = ({(operation_274_2619[7:0])});
    assign operation_274_2593 = ({(operation_274_2620[7:0])});
    assign operation_274_2592 = ({(operation_274_2621[7:0])});
    assign operation_274_2591 = ({(operation_274_2622[7:0])});
    assign operation_274_2589 = ({(operation_274_2623[7:0])});
    assign operation_274_2623 = (operation_274_2640);
    assign operation_274_2622 = (operation_274_2639);
    assign operation_274_2621 = (operation_274_2638);
    assign operation_274_2620 = (operation_274_2637);
    assign operation_274_2619 = (operation_274_2636);
    assign operation_274_2618 = (operation_274_2635);
    assign operation_274_2617 = (operation_274_2634);
    assign operation_274_2616 = (operation_274_2633);
    assign operation_274_2615 = (operation_274_2632);
    assign operation_274_2614 = (operation_274_2631);
    assign operation_274_2613 = (operation_274_2630);
    assign operation_274_2612 = (operation_274_2629);
    assign operation_274_2611 = (operation_274_2628);
    assign operation_274_2610 = (operation_274_2627);
    assign operation_274_2609 = (operation_274_2626);
    assign operation_274_2608 = (operation_274_2625);
    assign operation_274_3794 = ({(operation_274_3803[7:0])});
    assign operation_274_3793 = ({(operation_274_3804[7:0])});
    assign operation_274_3792 = ({(operation_274_3821[7:0])});
    assign operation_274_3775 = ({(operation_274_3822[7:0])});
    assign operation_274_3089 = ({(operation_274_3109[7:0])});
    assign operation_274_3088 = ({(operation_274_3108[7:0])});
    assign operation_274_3070 = ({(operation_274_3090[7:0])});
    assign operation_274_3019 = ({(operation_274_3036[7:0])});
    assign operation_274_3822 = ((control_274_23)?(lookup_sbox_0_output):(operation_274_3822_latch));
    assign operation_274_3821 = ((control_274_22)?(lookup_sbox_0_output):(operation_274_3821_latch));
    assign operation_274_3804 = ((control_274_22)?(lookup_sbox_1_output):(operation_274_3804_latch));
    assign operation_274_3803 = ((control_274_23)?(lookup_sbox_1_output):(operation_274_3803_latch));
    assign operation_274_2658 = ({(operation_274_2678[7:0])});
    assign operation_274_2657 = ({(operation_274_2677[7:0])});
    assign operation_274_2656 = ({(operation_274_2676[7:0])});
    assign operation_274_2655 = ({(operation_274_2675[7:0])});
    assign operation_274_2654 = ({(operation_274_2674[7:0])});
    assign operation_274_2653 = ({(operation_274_2673[7:0])});
    assign operation_274_2652 = ({(operation_274_2672[7:0])});
    assign operation_274_2651 = ({(operation_274_2671[7:0])});
    assign operation_274_2650 = ({(operation_274_2670[7:0])});
    assign operation_274_2649 = ({(operation_274_2669[7:0])});
    assign operation_274_2648 = ({(operation_274_2668[7:0])});
    assign operation_274_2647 = ({(operation_274_2667[7:0])});
    assign operation_274_2646 = ({(operation_274_2666[7:0])});
    assign operation_274_2645 = ({(operation_274_2665[7:0])});
    assign operation_274_2644 = ({(operation_274_2664[7:0])});
    assign operation_274_2643 = ({(operation_274_2663[7:0])});
    assign operation_274_3109 = (operation_274_3129);
    assign operation_274_3108 = (operation_274_3128);
    assign operation_274_3090 = (operation_274_3110);
    assign operation_274_3036 = (operation_274_3053);
    assign operation_274_2678 = (operation_274_2698);
    assign operation_274_2677 = (operation_274_2697);
    assign operation_274_2676 = (operation_274_2696);
    assign operation_274_2675 = (operation_274_2695);
    assign operation_274_2674 = (operation_274_2694);
    assign operation_274_2673 = (operation_274_2693);
    assign operation_274_2672 = (operation_274_2692);
    assign operation_274_2671 = (operation_274_2691);
    assign operation_274_2670 = (operation_274_2690);
    assign operation_274_2669 = (operation_274_2689);
    assign operation_274_2668 = (operation_274_2688);
    assign operation_274_2667 = (operation_274_2687);
    assign operation_274_2666 = (operation_274_2686);
    assign operation_274_2665 = (operation_274_2685);
    assign operation_274_2664 = (operation_274_2684);
    assign operation_274_2663 = (operation_274_2683);
    assign operation_274_3149 = ({(operation_274_3169[7:0])});
    assign operation_274_3148 = ({(operation_274_3168[7:0])});
    assign operation_274_3130 = ({(operation_274_3150[7:0])});
    assign operation_274_3071 = ({(operation_274_3091[7:0])});
    assign operation_274_2718 = ({(operation_274_2738[7:0])});
    assign operation_274_2717 = ({(operation_274_2737[7:0])});
    assign operation_274_2716 = ({(operation_274_2736[7:0])});
    assign operation_274_2715 = ({(operation_274_2735[7:0])});
    assign operation_274_2714 = ({(operation_274_2734[7:0])});
    assign operation_274_2713 = ({(operation_274_2733[7:0])});
    assign operation_274_2712 = ({(operation_274_2732[7:0])});
    assign operation_274_2711 = ({(operation_274_2731[7:0])});
    assign operation_274_2710 = ({(operation_274_2730[7:0])});
    assign operation_274_2709 = ({(operation_274_2729[7:0])});
    assign operation_274_2708 = ({(operation_274_2728[7:0])});
    assign operation_274_2707 = ({(operation_274_2727[7:0])});
    assign operation_274_2706 = ({(operation_274_2726[7:0])});
    assign operation_274_2705 = ({(operation_274_2725[7:0])});
    assign operation_274_2704 = ({(operation_274_2724[7:0])});
    assign operation_274_2703 = ({(operation_274_2723[7:0])});
    assign operation_274_3169 = (operation_274_3189);
    assign operation_274_3168 = (operation_274_3188);
    assign operation_274_3150 = (operation_274_3170);
    assign operation_274_3091 = (operation_274_3111);
    assign operation_274_2738 = (operation_274_2758);
    assign operation_274_2737 = (operation_274_2757);
    assign operation_274_2736 = (operation_274_2756);
    assign operation_274_2735 = (operation_274_2755);
    assign operation_274_2734 = (operation_274_2754);
    assign operation_274_2733 = (operation_274_2753);
    assign operation_274_2732 = (operation_274_2752);
    assign operation_274_2731 = (operation_274_2751);
    assign operation_274_2730 = (operation_274_2750);
    assign operation_274_2729 = (operation_274_2749);
    assign operation_274_2728 = (operation_274_2748);
    assign operation_274_2727 = (operation_274_2747);
    assign operation_274_2726 = (operation_274_2746);
    assign operation_274_2725 = (operation_274_2745);
    assign operation_274_2724 = (operation_274_2744);
    assign operation_274_2723 = (operation_274_2743);
    assign operation_274_3209 = ({(operation_274_3233[7:0])});
    assign operation_274_3208 = ({(operation_274_3232[7:0])});
    assign operation_274_3190 = ({(operation_274_3210[7:0])});
    assign operation_274_3131 = ({(operation_274_3151[7:0])});
    assign operation_274_3233 = (operation_274_3273);
    assign operation_274_3232 = (operation_274_3272);
    assign operation_274_3210 = (operation_274_3234);
    assign operation_274_3151 = (operation_274_3171);
    assign operation_274_2786 = ({(operation_274_2841[7:0])});
    assign operation_274_2785 = ({(operation_274_2808[7:0])});
    assign operation_274_2784 = ({(operation_274_2842[7:0])});
    assign operation_274_2783 = ({(operation_274_2807[7:0])});
    assign operation_274_2842 = (operation_274_2866);
    assign operation_274_2841 = (operation_274_2865);
    assign operation_274_2808 = (operation_274_2848);
    assign operation_274_2807 = (operation_274_2847);
    assign operation_274_3297 = ({(operation_274_3322[7:0])});
    assign operation_274_3296 = ({(operation_274_3321[7:0])});
    assign operation_274_3274 = ({(operation_274_3299[7:0])});
    assign operation_274_3191 = ({(operation_274_3211[7:0])});
    assign operation_274_2864 = ({(operation_274_2888[7:0])});
    assign operation_274_2863 = ({(operation_274_2887[7:0])});
    assign operation_274_2862 = ({(operation_274_2886[7:0])});
    assign operation_274_2861 = ({(operation_274_2885[7:0])});
    assign operation_274_2860 = ({(operation_274_2884[7:0])});
    assign operation_274_2859 = ({(operation_274_2883[7:0])});
    assign operation_274_2858 = ({(operation_274_2882[7:0])});
    assign operation_274_2857 = ({(operation_274_2881[7:0])});
    assign operation_274_2856 = ({(operation_274_2880[7:0])});
    assign operation_274_2855 = ({(operation_274_2879[7:0])});
    assign operation_274_2854 = ({(operation_274_2878[7:0])});
    assign operation_274_2853 = ({(operation_274_2877[7:0])});
    assign operation_274_2852 = ({(operation_274_2876[7:0])});
    assign operation_274_2851 = ({(operation_274_2875[7:0])});
    assign operation_274_2850 = ({(operation_274_2874[7:0])});
    assign operation_274_2849 = ({(operation_274_2873[7:0])});
    assign operation_274_3322 = (operation_274_3343);
    assign operation_274_3321 = (operation_274_3342);
    assign operation_274_3299 = (operation_274_3324);
    assign operation_274_3211 = (operation_274_3235);
    assign operation_274_2888 = (operation_274_2911);
    assign operation_274_2887 = (operation_274_2896);
    assign operation_274_2886 = (operation_274_2910);
    assign operation_274_2885 = (operation_274_2909);
    assign operation_274_2884 = (operation_274_2908);
    assign operation_274_2883 = (operation_274_2897);
    assign operation_274_2882 = (operation_274_2907);
    assign operation_274_2881 = (operation_274_2906);
    assign operation_274_2880 = (operation_274_2905);
    assign operation_274_2879 = (operation_274_2904);
    assign operation_274_2878 = (operation_274_2903);
    assign operation_274_2877 = (operation_274_2902);
    assign operation_274_2876 = (operation_274_2901);
    assign operation_274_2875 = (operation_274_2900);
    assign operation_274_2874 = (operation_274_2899);
    assign operation_274_2873 = (operation_274_2898);
    assign operation_274_3365 = ({(operation_274_3374[7:0])});
    assign operation_274_3364 = ({(operation_274_3375[7:0])});
    assign operation_274_3346 = ({(operation_274_3393[7:0])});
    assign operation_274_3275 = ({(operation_274_3320[7:0])});
    assign operation_274_2933 = ({(operation_274_2960[7:0])});
    assign operation_274_2932 = ({(operation_274_2955[7:0])});
    assign operation_274_2931 = ({(operation_274_2956[7:0])});
    assign operation_274_2930 = ({(operation_274_2959[7:0])});
    assign operation_274_2929 = ({(operation_274_2962[7:0])});
    assign operation_274_2928 = ({(operation_274_2957[7:0])});
    assign operation_274_2927 = ({(operation_274_2958[7:0])});
    assign operation_274_2926 = ({(operation_274_2961[7:0])});
    assign operation_274_2925 = ({(operation_274_2952[7:0])});
    assign operation_274_2924 = ({(operation_274_2947[7:0])});
    assign operation_274_2923 = ({(operation_274_2950[7:0])});
    assign operation_274_2922 = ({(operation_274_2953[7:0])});
    assign operation_274_2921 = ({(operation_274_2948[7:0])});
    assign operation_274_2920 = ({(operation_274_2951[7:0])});
    assign operation_274_2919 = ({(operation_274_2954[7:0])});
    assign operation_274_2918 = ({(operation_274_2949[7:0])});
    assign operation_274_2660 = ({(operation_274_2680[7:0])});
    assign operation_274_2641 = ({(operation_274_2661[7:0])});
    assign operation_274_2590 = ({(operation_274_2607[7:0])});
    assign operation_274_3393 = ((control_274_17)?(lookup_sbox_1_output):(operation_274_3393_latch));
    assign operation_274_3375 = ((control_274_17)?(lookup_sbox_2_output):(operation_274_3375_latch));
    assign operation_274_3374 = ((control_274_18)?(lookup_sbox_0_output):(operation_274_3374_latch));
    assign operation_274_3320 = (operation_274_3341);
    assign operation_274_2962 = ((control_274_20)?(lookup_sbox_0_output):(operation_274_2962_latch));
    assign operation_274_2961 = ((control_274_20)?(lookup_sbox_1_output):(operation_274_2961_latch));
    assign operation_274_2960 = ((control_274_20)?(lookup_sbox_2_output):(operation_274_2960_latch));
    assign operation_274_2959 = ((control_274_20)?(lookup_sbox_3_output):(operation_274_2959_latch));
    assign operation_274_2958 = ((control_274_20)?(lookup_sbox_4_output):(operation_274_2958_latch));
    assign operation_274_2957 = ((control_274_20)?(lookup_sbox_5_output):(operation_274_2957_latch));
    assign operation_274_2956 = ((control_274_20)?(lookup_sbox_6_output):(operation_274_2956_latch));
    assign operation_274_2955 = ((control_274_20)?(lookup_sbox_7_output):(operation_274_2955_latch));
    assign operation_274_2954 = ((control_274_20)?(lookup_sbox_8_output):(operation_274_2954_latch));
    assign operation_274_2953 = ((control_274_20)?(lookup_sbox_9_output):(operation_274_2953_latch));
    assign operation_274_2952 = ((control_274_20)?(lookup_sbox_10_output):(operation_274_2952_latch));
    assign operation_274_2951 = ((control_274_20)?(lookup_sbox_11_output):(operation_274_2951_latch));
    assign operation_274_2950 = ((control_274_20)?(lookup_sbox_12_output):(operation_274_2950_latch));
    assign operation_274_2949 = ((control_274_20)?(lookup_sbox_13_output):(operation_274_2949_latch));
    assign operation_274_2948 = ((control_274_20)?(lookup_sbox_14_output):(operation_274_2948_latch));
    assign operation_274_2947 = ((control_274_20)?(lookup_sbox_15_output):(operation_274_2947_latch));
    assign operation_274_2680 = (operation_274_2700);
    assign operation_274_2661 = (operation_274_2681);
    assign operation_274_2607 = (operation_274_2624);
    assign operation_274_2143 = (operation_274_2159);
    assign operation_274_2142 = (operation_274_2158);
    assign operation_274_2141 = (operation_274_2157);
    assign operation_274_2140 = (operation_274_2156);
    assign operation_274_2139 = (operation_274_2155);
    assign operation_274_2138 = (operation_274_2154);
    assign operation_274_2137 = (operation_274_2153);
    assign operation_274_2136 = (operation_274_2152);
    assign operation_274_2135 = (operation_274_2151);
    assign operation_274_2134 = (operation_274_2150);
    assign operation_274_2133 = (operation_274_2149);
    assign operation_274_2132 = (operation_274_2148);
    assign operation_274_2131 = (operation_274_2147);
    assign operation_274_2130 = (operation_274_2146);
    assign operation_274_2129 = (operation_274_2145);
    assign operation_274_2128 = (operation_274_2144);
    assign operation_274_3363 = ({(operation_274_3392[7:0])});
    assign operation_274_2720 = ({(operation_274_2740[7:0])});
    assign operation_274_2701 = ({(operation_274_2721[7:0])});
    assign operation_274_2659 = ({(operation_274_2679[7:0])});
    assign operation_274_2642 = ({(operation_274_2662[7:0])});
    assign operation_274_3392 = ((control_274_17)?(lookup_sbox_0_output):(operation_274_3392_latch));
    assign operation_274_2177 = ({(operation_274_2179[7:0])});
    assign operation_274_2176 = ({(operation_274_2180[7:0])});
    assign operation_274_2175 = ({(operation_274_2181[7:0])});
    assign operation_274_2174 = ({(operation_274_2182[7:0])});
    assign operation_274_2173 = ({(operation_274_2183[7:0])});
    assign operation_274_2172 = ({(operation_274_2184[7:0])});
    assign operation_274_2171 = ({(operation_274_2185[7:0])});
    assign operation_274_2170 = ({(operation_274_2186[7:0])});
    assign operation_274_2168 = ({(operation_274_2187[7:0])});
    assign operation_274_2167 = ({(operation_274_2188[7:0])});
    assign operation_274_2166 = ({(operation_274_2189[7:0])});
    assign operation_274_2165 = ({(operation_274_2190[7:0])});
    assign operation_274_2164 = ({(operation_274_2191[7:0])});
    assign operation_274_2163 = ({(operation_274_2192[7:0])});
    assign operation_274_2162 = ({(operation_274_2193[7:0])});
    assign operation_274_2160 = ({(operation_274_2194[7:0])});
    assign operation_274_2740 = (operation_274_2760);
    assign operation_274_2721 = (operation_274_2741);
    assign operation_274_2679 = (operation_274_2699);
    assign operation_274_2662 = (operation_274_2682);
    assign operation_274_2194 = (operation_274_2211);
    assign operation_274_2193 = (operation_274_2210);
    assign operation_274_2192 = (operation_274_2209);
    assign operation_274_2191 = (operation_274_2208);
    assign operation_274_2190 = (operation_274_2207);
    assign operation_274_2189 = (operation_274_2206);
    assign operation_274_2188 = (operation_274_2205);
    assign operation_274_2187 = (operation_274_2204);
    assign operation_274_2186 = (operation_274_2203);
    assign operation_274_2185 = (operation_274_2202);
    assign operation_274_2184 = (operation_274_2201);
    assign operation_274_2183 = (operation_274_2200);
    assign operation_274_2182 = (operation_274_2199);
    assign operation_274_2181 = (operation_274_2198);
    assign operation_274_2180 = (operation_274_2197);
    assign operation_274_2179 = (operation_274_2196);
    assign operation_274_2780 = ({(operation_274_2804[7:0])});
    assign operation_274_2761 = ({(operation_274_2781[7:0])});
    assign operation_274_2719 = ({(operation_274_2739[7:0])});
    assign operation_274_2702 = ({(operation_274_2722[7:0])});
    assign operation_274_2229 = ({(operation_274_2249[7:0])});
    assign operation_274_2228 = ({(operation_274_2248[7:0])});
    assign operation_274_2227 = ({(operation_274_2247[7:0])});
    assign operation_274_2226 = ({(operation_274_2246[7:0])});
    assign operation_274_2225 = ({(operation_274_2245[7:0])});
    assign operation_274_2224 = ({(operation_274_2244[7:0])});
    assign operation_274_2223 = ({(operation_274_2243[7:0])});
    assign operation_274_2222 = ({(operation_274_2242[7:0])});
    assign operation_274_2221 = ({(operation_274_2241[7:0])});
    assign operation_274_2220 = ({(operation_274_2240[7:0])});
    assign operation_274_2219 = ({(operation_274_2239[7:0])});
    assign operation_274_2218 = ({(operation_274_2238[7:0])});
    assign operation_274_2217 = ({(operation_274_2237[7:0])});
    assign operation_274_2216 = ({(operation_274_2236[7:0])});
    assign operation_274_2215 = ({(operation_274_2235[7:0])});
    assign operation_274_2214 = ({(operation_274_2234[7:0])});
    assign operation_274_2804 = (operation_274_2844);
    assign operation_274_2781 = (operation_274_2805);
    assign operation_274_2739 = (operation_274_2759);
    assign operation_274_2722 = (operation_274_2742);
    assign operation_274_2249 = (operation_274_2269);
    assign operation_274_2248 = (operation_274_2268);
    assign operation_274_2247 = (operation_274_2267);
    assign operation_274_2246 = (operation_274_2266);
    assign operation_274_2245 = (operation_274_2265);
    assign operation_274_2244 = (operation_274_2264);
    assign operation_274_2243 = (operation_274_2263);
    assign operation_274_2242 = (operation_274_2262);
    assign operation_274_2241 = (operation_274_2261);
    assign operation_274_2240 = (operation_274_2260);
    assign operation_274_2239 = (operation_274_2259);
    assign operation_274_2238 = (operation_274_2258);
    assign operation_274_2237 = (operation_274_2257);
    assign operation_274_2236 = (operation_274_2256);
    assign operation_274_2235 = (operation_274_2255);
    assign operation_274_2234 = (operation_274_2254);
    assign operation_274_2868 = ({(operation_274_2893[7:0])});
    assign operation_274_2845 = ({(operation_274_2870[7:0])});
    assign operation_274_2779 = ({(operation_274_2803[7:0])});
    assign operation_274_2762 = ({(operation_274_2782[7:0])});
    assign operation_274_2289 = ({(operation_274_2309[7:0])});
    assign operation_274_2288 = ({(operation_274_2308[7:0])});
    assign operation_274_2287 = ({(operation_274_2307[7:0])});
    assign operation_274_2286 = ({(operation_274_2306[7:0])});
    assign operation_274_2285 = ({(operation_274_2305[7:0])});
    assign operation_274_2284 = ({(operation_274_2304[7:0])});
    assign operation_274_2283 = ({(operation_274_2303[7:0])});
    assign operation_274_2282 = ({(operation_274_2302[7:0])});
    assign operation_274_2281 = ({(operation_274_2301[7:0])});
    assign operation_274_2280 = ({(operation_274_2300[7:0])});
    assign operation_274_2279 = ({(operation_274_2299[7:0])});
    assign operation_274_2278 = ({(operation_274_2298[7:0])});
    assign operation_274_2277 = ({(operation_274_2297[7:0])});
    assign operation_274_2276 = ({(operation_274_2296[7:0])});
    assign operation_274_2275 = ({(operation_274_2295[7:0])});
    assign operation_274_2274 = ({(operation_274_2294[7:0])});
    assign operation_274_2893 = (operation_274_2914);
    assign operation_274_2870 = (operation_274_2895);
    assign operation_274_2803 = (operation_274_2843);
    assign operation_274_2782 = (operation_274_2806);
    assign operation_274_2309 = (operation_274_2329);
    assign operation_274_2308 = (operation_274_2328);
    assign operation_274_2307 = (operation_274_2327);
    assign operation_274_2306 = (operation_274_2326);
    assign operation_274_2305 = (operation_274_2325);
    assign operation_274_2304 = (operation_274_2324);
    assign operation_274_2303 = (operation_274_2323);
    assign operation_274_2302 = (operation_274_2322);
    assign operation_274_2301 = (operation_274_2321);
    assign operation_274_2300 = (operation_274_2320);
    assign operation_274_2299 = (operation_274_2319);
    assign operation_274_2298 = (operation_274_2318);
    assign operation_274_2297 = (operation_274_2317);
    assign operation_274_2296 = (operation_274_2316);
    assign operation_274_2295 = (operation_274_2315);
    assign operation_274_2294 = (operation_274_2314);
    assign operation_274_2936 = ({(operation_274_2945[7:0])});
    assign operation_274_2917 = ({(operation_274_2964[7:0])});
    assign operation_274_2867 = ({(operation_274_2892[7:0])});
    assign operation_274_2846 = ({(operation_274_2891[7:0])});
    assign operation_274_2231 = ({(operation_274_2251[7:0])});
    assign operation_274_2161 = ({(operation_274_2178[7:0])});
    assign operation_274_2964 = ((control_274_12)?(lookup_sbox_2_output):(operation_274_2964_latch));
    assign operation_274_2945 = ((control_274_12)?(lookup_sbox_3_output):(operation_274_2945_latch));
    assign operation_274_2892 = (operation_274_2913);
    assign operation_274_2891 = (operation_274_2912);
    assign operation_274_2357 = ({(operation_274_2412[7:0])});
    assign operation_274_2356 = ({(operation_274_2379[7:0])});
    assign operation_274_2355 = ({(operation_274_2413[7:0])});
    assign operation_274_2354 = ({(operation_274_2378[7:0])});
    assign operation_274_2251 = (operation_274_2271);
    assign operation_274_2178 = (operation_274_2195);
    assign operation_274_2413 = (operation_274_2437);
    assign operation_274_2412 = (operation_274_2436);
    assign operation_274_2379 = (operation_274_2419);
    assign operation_274_2378 = (operation_274_2418);
    assign operation_274_2935 = ({(operation_274_2946[7:0])});
    assign operation_274_2934 = ({(operation_274_2963[7:0])});
    assign operation_274_2435 = ({(operation_274_2459[7:0])});
    assign operation_274_2434 = ({(operation_274_2458[7:0])});
    assign operation_274_2433 = ({(operation_274_2457[7:0])});
    assign operation_274_2432 = ({(operation_274_2456[7:0])});
    assign operation_274_2431 = ({(operation_274_2455[7:0])});
    assign operation_274_2430 = ({(operation_274_2454[7:0])});
    assign operation_274_2429 = ({(operation_274_2453[7:0])});
    assign operation_274_2428 = ({(operation_274_2452[7:0])});
    assign operation_274_2427 = ({(operation_274_2451[7:0])});
    assign operation_274_2426 = ({(operation_274_2450[7:0])});
    assign operation_274_2425 = ({(operation_274_2449[7:0])});
    assign operation_274_2424 = ({(operation_274_2448[7:0])});
    assign operation_274_2423 = ({(operation_274_2447[7:0])});
    assign operation_274_2422 = ({(operation_274_2446[7:0])});
    assign operation_274_2421 = ({(operation_274_2445[7:0])});
    assign operation_274_2420 = ({(operation_274_2444[7:0])});
    assign operation_274_2291 = ({(operation_274_2311[7:0])});
    assign operation_274_2230 = ({(operation_274_2250[7:0])});
    assign operation_274_2213 = ({(operation_274_2233[7:0])});
    assign operation_274_2212 = ({(operation_274_2232[7:0])});
    assign operation_274_2963 = ((control_274_12)?(lookup_sbox_0_output):(operation_274_2963_latch));
    assign operation_274_2946 = ((control_274_12)?(lookup_sbox_1_output):(operation_274_2946_latch));
    assign operation_274_2459 = (operation_274_2482);
    assign operation_274_2458 = (operation_274_2467);
    assign operation_274_2457 = (operation_274_2481);
    assign operation_274_2456 = (operation_274_2480);
    assign operation_274_2455 = (operation_274_2479);
    assign operation_274_2454 = (operation_274_2468);
    assign operation_274_2453 = (operation_274_2478);
    assign operation_274_2452 = (operation_274_2477);
    assign operation_274_2451 = (operation_274_2476);
    assign operation_274_2450 = (operation_274_2475);
    assign operation_274_2449 = (operation_274_2474);
    assign operation_274_2448 = (operation_274_2473);
    assign operation_274_2447 = (operation_274_2472);
    assign operation_274_2446 = (operation_274_2471);
    assign operation_274_2445 = (operation_274_2470);
    assign operation_274_2444 = (operation_274_2469);
    assign operation_274_2311 = (operation_274_2331);
    assign operation_274_2250 = (operation_274_2270);
    assign operation_274_2233 = (operation_274_2253);
    assign operation_274_2232 = (operation_274_2252);
    assign operation_274_2504 = ({(operation_274_2531[7:0])});
    assign operation_274_2503 = ({(operation_274_2526[7:0])});
    assign operation_274_2502 = ({(operation_274_2527[7:0])});
    assign operation_274_2501 = ({(operation_274_2530[7:0])});
    assign operation_274_2500 = ({(operation_274_2533[7:0])});
    assign operation_274_2499 = ({(operation_274_2528[7:0])});
    assign operation_274_2498 = ({(operation_274_2529[7:0])});
    assign operation_274_2497 = ({(operation_274_2532[7:0])});
    assign operation_274_2496 = ({(operation_274_2523[7:0])});
    assign operation_274_2495 = ({(operation_274_2518[7:0])});
    assign operation_274_2494 = ({(operation_274_2521[7:0])});
    assign operation_274_2493 = ({(operation_274_2524[7:0])});
    assign operation_274_2492 = ({(operation_274_2519[7:0])});
    assign operation_274_2491 = ({(operation_274_2522[7:0])});
    assign operation_274_2490 = ({(operation_274_2525[7:0])});
    assign operation_274_2489 = ({(operation_274_2520[7:0])});
    assign operation_274_2351 = ({(operation_274_2375[7:0])});
    assign operation_274_2290 = ({(operation_274_2310[7:0])});
    assign operation_274_2273 = ({(operation_274_2293[7:0])});
    assign operation_274_2272 = ({(operation_274_2292[7:0])});
    assign operation_274_2533 = ((control_274_11)?(lookup_sbox_0_output):(operation_274_2533_latch));
    assign operation_274_2532 = ((control_274_11)?(lookup_sbox_1_output):(operation_274_2532_latch));
    assign operation_274_2531 = ((control_274_11)?(lookup_sbox_2_output):(operation_274_2531_latch));
    assign operation_274_2530 = ((control_274_11)?(lookup_sbox_3_output):(operation_274_2530_latch));
    assign operation_274_2529 = ((control_274_11)?(lookup_sbox_4_output):(operation_274_2529_latch));
    assign operation_274_2528 = ((control_274_11)?(lookup_sbox_5_output):(operation_274_2528_latch));
    assign operation_274_2527 = ((control_274_11)?(lookup_sbox_6_output):(operation_274_2527_latch));
    assign operation_274_2526 = ((control_274_11)?(lookup_sbox_7_output):(operation_274_2526_latch));
    assign operation_274_2525 = ((control_274_11)?(lookup_sbox_8_output):(operation_274_2525_latch));
    assign operation_274_2524 = ((control_274_11)?(lookup_sbox_9_output):(operation_274_2524_latch));
    assign operation_274_2523 = ((control_274_11)?(lookup_sbox_10_output):(operation_274_2523_latch));
    assign operation_274_2522 = ((control_274_11)?(lookup_sbox_11_output):(operation_274_2522_latch));
    assign operation_274_2521 = ((control_274_11)?(lookup_sbox_12_output):(operation_274_2521_latch));
    assign operation_274_2520 = ((control_274_11)?(lookup_sbox_13_output):(operation_274_2520_latch));
    assign operation_274_2519 = ((control_274_11)?(lookup_sbox_14_output):(operation_274_2519_latch));
    assign operation_274_2518 = ((control_274_11)?(lookup_sbox_15_output):(operation_274_2518_latch));
    assign operation_274_2375 = (operation_274_2415);
    assign operation_274_2310 = (operation_274_2330);
    assign operation_274_2293 = (operation_274_2313);
    assign operation_274_2292 = (operation_274_2312);
    assign operation_274_1714 = (operation_274_1730);
    assign operation_274_1713 = (operation_274_1729);
    assign operation_274_1712 = (operation_274_1728);
    assign operation_274_1711 = (operation_274_1727);
    assign operation_274_1710 = (operation_274_1726);
    assign operation_274_1709 = (operation_274_1725);
    assign operation_274_1708 = (operation_274_1724);
    assign operation_274_1707 = (operation_274_1723);
    assign operation_274_1706 = (operation_274_1722);
    assign operation_274_1705 = (operation_274_1721);
    assign operation_274_1704 = (operation_274_1720);
    assign operation_274_1703 = (operation_274_1719);
    assign operation_274_1702 = (operation_274_1718);
    assign operation_274_1701 = (operation_274_1717);
    assign operation_274_1700 = (operation_274_1716);
    assign operation_274_1699 = (operation_274_1715);
    assign operation_274_2439 = ({(operation_274_2464[7:0])});
    assign operation_274_2350 = ({(operation_274_2374[7:0])});
    assign operation_274_2333 = ({(operation_274_2353[7:0])});
    assign operation_274_2332 = ({(operation_274_2352[7:0])});
    assign operation_274_1748 = ({(operation_274_1750[7:0])});
    assign operation_274_1747 = ({(operation_274_1751[7:0])});
    assign operation_274_1746 = ({(operation_274_1752[7:0])});
    assign operation_274_1745 = ({(operation_274_1753[7:0])});
    assign operation_274_1744 = ({(operation_274_1754[7:0])});
    assign operation_274_1743 = ({(operation_274_1755[7:0])});
    assign operation_274_1742 = ({(operation_274_1756[7:0])});
    assign operation_274_1741 = ({(operation_274_1757[7:0])});
    assign operation_274_1739 = ({(operation_274_1758[7:0])});
    assign operation_274_1738 = ({(operation_274_1759[7:0])});
    assign operation_274_1737 = ({(operation_274_1760[7:0])});
    assign operation_274_1736 = ({(operation_274_1761[7:0])});
    assign operation_274_1735 = ({(operation_274_1762[7:0])});
    assign operation_274_1734 = ({(operation_274_1763[7:0])});
    assign operation_274_1733 = ({(operation_274_1764[7:0])});
    assign operation_274_1731 = ({(operation_274_1765[7:0])});
    assign operation_274_2464 = (operation_274_2485);
    assign operation_274_2374 = (operation_274_2414);
    assign operation_274_2353 = (operation_274_2377);
    assign operation_274_2352 = (operation_274_2376);
    assign operation_274_1765 = (operation_274_1782);
    assign operation_274_1764 = (operation_274_1781);
    assign operation_274_1763 = (operation_274_1780);
    assign operation_274_1762 = (operation_274_1779);
    assign operation_274_1761 = (operation_274_1778);
    assign operation_274_1760 = (operation_274_1777);
    assign operation_274_1759 = (operation_274_1776);
    assign operation_274_1758 = (operation_274_1775);
    assign operation_274_1757 = (operation_274_1774);
    assign operation_274_1756 = (operation_274_1773);
    assign operation_274_1755 = (operation_274_1772);
    assign operation_274_1754 = (operation_274_1771);
    assign operation_274_1753 = (operation_274_1770);
    assign operation_274_1752 = (operation_274_1769);
    assign operation_274_1751 = (operation_274_1768);
    assign operation_274_1750 = (operation_274_1767);
    assign operation_274_2507 = ({(operation_274_2516[7:0])});
    assign operation_274_2438 = ({(operation_274_2463[7:0])});
    assign operation_274_2417 = ({(operation_274_2462[7:0])});
    assign operation_274_2416 = ({(operation_274_2441[7:0])});
    assign operation_274_1800 = ({(operation_274_1820[7:0])});
    assign operation_274_1799 = ({(operation_274_1819[7:0])});
    assign operation_274_1798 = ({(operation_274_1818[7:0])});
    assign operation_274_1797 = ({(operation_274_1817[7:0])});
    assign operation_274_1796 = ({(operation_274_1816[7:0])});
    assign operation_274_1795 = ({(operation_274_1815[7:0])});
    assign operation_274_1794 = ({(operation_274_1814[7:0])});
    assign operation_274_1793 = ({(operation_274_1813[7:0])});
    assign operation_274_1792 = ({(operation_274_1812[7:0])});
    assign operation_274_1791 = ({(operation_274_1811[7:0])});
    assign operation_274_1790 = ({(operation_274_1810[7:0])});
    assign operation_274_1789 = ({(operation_274_1809[7:0])});
    assign operation_274_1788 = ({(operation_274_1808[7:0])});
    assign operation_274_1787 = ({(operation_274_1807[7:0])});
    assign operation_274_1786 = ({(operation_274_1806[7:0])});
    assign operation_274_1785 = ({(operation_274_1805[7:0])});
    assign operation_274_1732 = ({(operation_274_1749[7:0])});
    assign operation_274_2516 = ((control_274_7)?(lookup_sbox_0_output):(operation_274_2516_latch));
    assign operation_274_2463 = (operation_274_2484);
    assign operation_274_2462 = (operation_274_2483);
    assign operation_274_2441 = (operation_274_2466);
    assign operation_274_1820 = (operation_274_1840);
    assign operation_274_1819 = (operation_274_1839);
    assign operation_274_1818 = (operation_274_1838);
    assign operation_274_1817 = (operation_274_1837);
    assign operation_274_1816 = (operation_274_1836);
    assign operation_274_1815 = (operation_274_1835);
    assign operation_274_1814 = (operation_274_1834);
    assign operation_274_1813 = (operation_274_1833);
    assign operation_274_1812 = (operation_274_1832);
    assign operation_274_1811 = (operation_274_1831);
    assign operation_274_1810 = (operation_274_1830);
    assign operation_274_1809 = (operation_274_1829);
    assign operation_274_1808 = (operation_274_1828);
    assign operation_274_1807 = (operation_274_1827);
    assign operation_274_1806 = (operation_274_1826);
    assign operation_274_1805 = (operation_274_1825);
    assign operation_274_1749 = (operation_274_1766);
    assign operation_274_2506 = ({(operation_274_2517[7:0])});
    assign operation_274_2505 = ({(operation_274_2534[7:0])});
    assign operation_274_2488 = ({(operation_274_2535[7:0])});
    assign operation_274_1860 = ({(operation_274_1880[7:0])});
    assign operation_274_1859 = ({(operation_274_1879[7:0])});
    assign operation_274_1858 = ({(operation_274_1878[7:0])});
    assign operation_274_1857 = ({(operation_274_1877[7:0])});
    assign operation_274_1856 = ({(operation_274_1876[7:0])});
    assign operation_274_1855 = ({(operation_274_1875[7:0])});
    assign operation_274_1854 = ({(operation_274_1874[7:0])});
    assign operation_274_1853 = ({(operation_274_1873[7:0])});
    assign operation_274_1852 = ({(operation_274_1872[7:0])});
    assign operation_274_1851 = ({(operation_274_1871[7:0])});
    assign operation_274_1850 = ({(operation_274_1870[7:0])});
    assign operation_274_1849 = ({(operation_274_1869[7:0])});
    assign operation_274_1848 = ({(operation_274_1868[7:0])});
    assign operation_274_1847 = ({(operation_274_1867[7:0])});
    assign operation_274_1846 = ({(operation_274_1866[7:0])});
    assign operation_274_1845 = ({(operation_274_1865[7:0])});
    assign operation_274_1802 = ({(operation_274_1822[7:0])});
    assign operation_274_1801 = ({(operation_274_1821[7:0])});
    assign operation_274_1784 = ({(operation_274_1804[7:0])});
    assign operation_274_1783 = ({(operation_274_1803[7:0])});
    assign operation_274_2535 = ((control_274_6)?(lookup_sbox_1_output):(operation_274_2535_latch));
    assign operation_274_2534 = ((control_274_6)?(lookup_sbox_0_output):(operation_274_2534_latch));
    assign operation_274_2517 = ((control_274_6)?(lookup_sbox_2_output):(operation_274_2517_latch));
    assign operation_274_1880 = (operation_274_1900);
    assign operation_274_1879 = (operation_274_1899);
    assign operation_274_1878 = (operation_274_1898);
    assign operation_274_1877 = (operation_274_1897);
    assign operation_274_1876 = (operation_274_1896);
    assign operation_274_1875 = (operation_274_1895);
    assign operation_274_1874 = (operation_274_1894);
    assign operation_274_1873 = (operation_274_1893);
    assign operation_274_1872 = (operation_274_1892);
    assign operation_274_1871 = (operation_274_1891);
    assign operation_274_1870 = (operation_274_1890);
    assign operation_274_1869 = (operation_274_1889);
    assign operation_274_1868 = (operation_274_1888);
    assign operation_274_1867 = (operation_274_1887);
    assign operation_274_1866 = (operation_274_1886);
    assign operation_274_1865 = (operation_274_1885);
    assign operation_274_1822 = (operation_274_1842);
    assign operation_274_1821 = (operation_274_1841);
    assign operation_274_1804 = (operation_274_1824);
    assign operation_274_1803 = (operation_274_1823);
    assign operation_274_1862 = ({(operation_274_1882[7:0])});
    assign operation_274_1861 = ({(operation_274_1881[7:0])});
    assign operation_274_1844 = ({(operation_274_1864[7:0])});
    assign operation_274_1843 = ({(operation_274_1863[7:0])});
    assign operation_274_1928 = ({(operation_274_1983[7:0])});
    assign operation_274_1927 = ({(operation_274_1950[7:0])});
    assign operation_274_1926 = ({(operation_274_1984[7:0])});
    assign operation_274_1925 = ({(operation_274_1949[7:0])});
    assign operation_274_1882 = (operation_274_1902);
    assign operation_274_1881 = (operation_274_1901);
    assign operation_274_1864 = (operation_274_1884);
    assign operation_274_1863 = (operation_274_1883);
    assign operation_274_1984 = (operation_274_2008);
    assign operation_274_1983 = (operation_274_2007);
    assign operation_274_1950 = (operation_274_1990);
    assign operation_274_1949 = (operation_274_1989);
    assign operation_274_2006 = ({(operation_274_2030[7:0])});
    assign operation_274_2005 = ({(operation_274_2029[7:0])});
    assign operation_274_2004 = ({(operation_274_2028[7:0])});
    assign operation_274_2003 = ({(operation_274_2027[7:0])});
    assign operation_274_2002 = ({(operation_274_2026[7:0])});
    assign operation_274_2001 = ({(operation_274_2025[7:0])});
    assign operation_274_2000 = ({(operation_274_2024[7:0])});
    assign operation_274_1999 = ({(operation_274_2023[7:0])});
    assign operation_274_1998 = ({(operation_274_2022[7:0])});
    assign operation_274_1997 = ({(operation_274_2021[7:0])});
    assign operation_274_1996 = ({(operation_274_2020[7:0])});
    assign operation_274_1995 = ({(operation_274_2019[7:0])});
    assign operation_274_1994 = ({(operation_274_2018[7:0])});
    assign operation_274_1993 = ({(operation_274_2017[7:0])});
    assign operation_274_1992 = ({(operation_274_2016[7:0])});
    assign operation_274_1991 = ({(operation_274_2015[7:0])});
    assign operation_274_1922 = ({(operation_274_1946[7:0])});
    assign operation_274_1921 = ({(operation_274_1945[7:0])});
    assign operation_274_1904 = ({(operation_274_1924[7:0])});
    assign operation_274_1903 = ({(operation_274_1923[7:0])});
    assign operation_274_2030 = (operation_274_2053);
    assign operation_274_2029 = (operation_274_2038);
    assign operation_274_2028 = (operation_274_2052);
    assign operation_274_2027 = (operation_274_2051);
    assign operation_274_2026 = (operation_274_2050);
    assign operation_274_2025 = (operation_274_2039);
    assign operation_274_2024 = (operation_274_2049);
    assign operation_274_2023 = (operation_274_2048);
    assign operation_274_2022 = (operation_274_2047);
    assign operation_274_2021 = (operation_274_2046);
    assign operation_274_2020 = (operation_274_2045);
    assign operation_274_2019 = (operation_274_2044);
    assign operation_274_2018 = (operation_274_2043);
    assign operation_274_2017 = (operation_274_2042);
    assign operation_274_2016 = (operation_274_2041);
    assign operation_274_2015 = (operation_274_2040);
    assign operation_274_1946 = (operation_274_1986);
    assign operation_274_1945 = (operation_274_1985);
    assign operation_274_1924 = (operation_274_1948);
    assign operation_274_1923 = (operation_274_1947);
    assign operation_274_2075 = ({(operation_274_2102[7:0])});
    assign operation_274_2074 = ({(operation_274_2097[7:0])});
    assign operation_274_2073 = ({(operation_274_2098[7:0])});
    assign operation_274_2072 = ({(operation_274_2101[7:0])});
    assign operation_274_2071 = ({(operation_274_2104[7:0])});
    assign operation_274_2070 = ({(operation_274_2099[7:0])});
    assign operation_274_2069 = ({(operation_274_2100[7:0])});
    assign operation_274_2068 = ({(operation_274_2103[7:0])});
    assign operation_274_2067 = ({(operation_274_2094[7:0])});
    assign operation_274_2066 = ({(operation_274_2089[7:0])});
    assign operation_274_2065 = ({(operation_274_2092[7:0])});
    assign operation_274_2064 = ({(operation_274_2095[7:0])});
    assign operation_274_2063 = ({(operation_274_2090[7:0])});
    assign operation_274_2062 = ({(operation_274_2093[7:0])});
    assign operation_274_2061 = ({(operation_274_2096[7:0])});
    assign operation_274_2060 = ({(operation_274_2091[7:0])});
    assign operation_274_2010 = ({(operation_274_2035[7:0])});
    assign operation_274_2009 = ({(operation_274_2034[7:0])});
    assign operation_274_1988 = ({(operation_274_2033[7:0])});
    assign operation_274_1987 = ({(operation_274_2012[7:0])});
    assign operation_274_2104 = ((control_274_2)?(lookup_sbox_0_output):(operation_274_2104_latch));
    assign operation_274_2103 = ((control_274_2)?(lookup_sbox_1_output):(operation_274_2103_latch));
    assign operation_274_2102 = ((control_274_2)?(lookup_sbox_2_output):(operation_274_2102_latch));
    assign operation_274_2101 = ((control_274_2)?(lookup_sbox_3_output):(operation_274_2101_latch));
    assign operation_274_2100 = ((control_274_2)?(lookup_sbox_4_output):(operation_274_2100_latch));
    assign operation_274_2099 = ((control_274_2)?(lookup_sbox_5_output):(operation_274_2099_latch));
    assign operation_274_2098 = ((control_274_2)?(lookup_sbox_6_output):(operation_274_2098_latch));
    assign operation_274_2097 = ((control_274_2)?(lookup_sbox_7_output):(operation_274_2097_latch));
    assign operation_274_2096 = ((control_274_2)?(lookup_sbox_8_output):(operation_274_2096_latch));
    assign operation_274_2095 = ((control_274_2)?(lookup_sbox_9_output):(operation_274_2095_latch));
    assign operation_274_2094 = ((control_274_2)?(lookup_sbox_10_output):(operation_274_2094_latch));
    assign operation_274_2093 = ((control_274_2)?(lookup_sbox_11_output):(operation_274_2093_latch));
    assign operation_274_2092 = ((control_274_2)?(lookup_sbox_12_output):(operation_274_2092_latch));
    assign operation_274_2091 = ((control_274_2)?(lookup_sbox_13_output):(operation_274_2091_latch));
    assign operation_274_2090 = ((control_274_2)?(lookup_sbox_14_output):(operation_274_2090_latch));
    assign operation_274_2089 = ((control_274_2)?(lookup_sbox_15_output):(operation_274_2089_latch));
    assign operation_274_2035 = (operation_274_2056);
    assign operation_274_2034 = (operation_274_2055);
    assign operation_274_2033 = (operation_274_2054);
    assign operation_274_2012 = (operation_274_2037);
    assign operation_274_119 = (operation_274_118);
    assign operation_274_103 = (operation_274_102);
    assign operation_274_87 = (operation_274_86);
    assign operation_274_71 = (operation_274_70);
    assign operation_274_55 = (operation_274_54);
    assign operation_274_39 = (operation_274_38);
    assign operation_274_23 = (operation_274_22);
    assign operation_274_7 = (operation_274_6);
    assign operation_274_15 = (operation_274_14);
    assign operation_274_31 = (operation_274_30);
    assign operation_274_47 = (operation_274_46);
    assign operation_274_63 = (operation_274_62);
    assign operation_274_79 = (operation_274_78);
    assign operation_274_95 = (operation_274_94);
    assign operation_274_111 = (operation_274_110);
    assign operation_274_127 = (operation_274_126);
    assign operation_274_2078 = ({(operation_274_2087[7:0])});
    assign operation_274_2077 = ({(operation_274_2088[7:0])});
    assign operation_274_2076 = ({(operation_274_2105[7:0])});
    assign operation_274_2059 = ({(operation_274_2106[7:0])});
    assign operation_274_117 = ({(operation_274_124[119:112])});
    assign operation_274_115 = ({(operation_274_122[119:112])});
    assign operation_274_101 = ({(operation_274_124[103:96])});
    assign operation_274_99 = ({(operation_274_122[103:96])});
    assign operation_274_85 = ({(operation_274_124[87:80])});
    assign operation_274_83 = ({(operation_274_122[87:80])});
    assign operation_274_69 = ({(operation_274_124[71:64])});
    assign operation_274_67 = ({(operation_274_122[71:64])});
    assign operation_274_53 = ({(operation_274_124[55:48])});
    assign operation_274_51 = ({(operation_274_122[55:48])});
    assign operation_274_37 = ({(operation_274_124[39:32])});
    assign operation_274_35 = ({(operation_274_122[39:32])});
    assign operation_274_21 = ({(operation_274_124[23:16])});
    assign operation_274_19 = ({(operation_274_122[23:16])});
    assign operation_274_5 = ({(operation_274_124[7:0])});
    assign operation_274_3 = ({(operation_274_122[7:0])});
    assign operation_274_11 = ({(operation_274_122[15:8])});
    assign operation_274_13 = ({(operation_274_124[15:8])});
    assign operation_274_27 = ({(operation_274_122[31:24])});
    assign operation_274_29 = ({(operation_274_124[31:24])});
    assign operation_274_43 = ({(operation_274_122[47:40])});
    assign operation_274_45 = ({(operation_274_124[47:40])});
    assign operation_274_59 = ({(operation_274_122[63:56])});
    assign operation_274_61 = ({(operation_274_124[63:56])});
    assign operation_274_75 = ({(operation_274_122[79:72])});
    assign operation_274_77 = ({(operation_274_124[79:72])});
    assign operation_274_91 = ({(operation_274_122[95:88])});
    assign operation_274_93 = ({(operation_274_124[95:88])});
    assign operation_274_107 = ({(operation_274_122[111:104])});
    assign operation_274_109 = ({(operation_274_124[111:104])});
    assign operation_274_123 = ({(operation_274_122[127:120])});
    assign operation_274_125 = ({(operation_274_124[127:120])});
    assign operation_274_2106 = ((control_274_1)?(lookup_sbox_1_output):(operation_274_2106_latch));
    assign operation_274_2105 = ((control_274_1)?(lookup_sbox_0_output):(operation_274_2105_latch));
    assign operation_274_2088 = ((control_274_1)?(lookup_sbox_2_output):(operation_274_2088_latch));
    assign operation_274_2087 = ((control_274_1)?(lookup_sbox_3_output):(operation_274_2087_latch));
    assign operation_274_5601 = (32'd54);
    assign operation_274_5597 = (32'd27);
    assign operation_274_5592 = (32'd128);
    assign operation_274_5587 = (32'd64);
    assign operation_274_5582 = (32'd32);
    assign operation_274_5577 = (32'd16);
    assign operation_274_5572 = (32'd8);
    assign operation_274_5567 = (32'd4);
    assign operation_274_5562 = (32'd2);
    assign operation_274_5557 = (32'd1);
    assign operation_274_2119 = (32'd7);
    assign operation_274_124 = (input_key_274);
    assign operation_274_122 = (input_in_274);
    assign control_274_end = (control_274_84);
    assign control_274_0 = (control_274_start);
    
    always_ff @(posedge clk)
    if(rst)
         begin
            finish <= 1'd0;
            AES128_encrypt <= 128'd0;
            operation_274_1664 <= 32'd0;
            operation_274_1688 <= 32'd0;
            operation_274_1672 <= 32'd0;
            operation_274_1632 <= 32'd0;
            operation_274_1680 <= 32'd0;
            operation_274_1656 <= 32'd0;
            operation_274_1640 <= 32'd0;
            operation_274_1600 <= 32'd0;
            operation_274_1648 <= 32'd0;
            operation_274_1624 <= 32'd0;
            operation_274_1608 <= 32'd0;
            operation_274_1568 <= 32'd0;
            operation_274_1616 <= 32'd0;
            operation_274_1592 <= 32'd0;
            operation_274_1576 <= 32'd0;
            operation_274_1584 <= 32'd0;
            operation_274_1338_latch <= 8'd0;
            operation_274_1328_latch <= 8'd0;
            operation_274_1318_latch <= 8'd0;
            operation_274_1308_latch <= 8'd0;
            operation_274_1298_latch <= 8'd0;
            operation_274_1288_latch <= 8'd0;
            operation_274_1278_latch <= 8'd0;
            operation_274_1268_latch <= 8'd0;
            operation_274_1273_latch <= 8'd0;
            operation_274_1283_latch <= 8'd0;
            operation_274_1293_latch <= 8'd0;
            operation_274_1303_latch <= 8'd0;
            operation_274_1313_latch <= 8'd0;
            operation_274_1323_latch <= 8'd0;
            operation_274_1333_latch <= 8'd0;
            operation_274_1343_latch <= 8'd0;
            operation_274_5162 <= 32'd0;
            operation_274_5161 <= 32'd0;
            operation_274_5160 <= 32'd0;
            operation_274_5159 <= 32'd0;
            operation_274_5158 <= 32'd0;
            operation_274_5157 <= 32'd0;
            operation_274_5156 <= 32'd0;
            operation_274_5155 <= 32'd0;
            operation_274_5154 <= 32'd0;
            operation_274_5153 <= 32'd0;
            operation_274_5152 <= 32'd0;
            operation_274_5151 <= 32'd0;
            operation_274_5150 <= 32'd0;
            operation_274_5149 <= 32'd0;
            operation_274_5148 <= 32'd0;
            operation_274_5147 <= 32'd0;
            operation_274_5214 <= 32'd0;
            operation_274_5213 <= 32'd0;
            operation_274_5212 <= 32'd0;
            operation_274_5211 <= 32'd0;
            operation_274_5210 <= 32'd0;
            operation_274_5209 <= 32'd0;
            operation_274_5208 <= 32'd0;
            operation_274_5207 <= 32'd0;
            operation_274_5206 <= 32'd0;
            operation_274_5205 <= 32'd0;
            operation_274_5204 <= 32'd0;
            operation_274_5203 <= 32'd0;
            operation_274_5202 <= 32'd0;
            operation_274_5201 <= 32'd0;
            operation_274_5200 <= 32'd0;
            operation_274_5199 <= 32'd0;
            operation_274_5272 <= 32'd0;
            operation_274_5271 <= 32'd0;
            operation_274_5270 <= 32'd0;
            operation_274_5269 <= 32'd0;
            operation_274_5268 <= 32'd0;
            operation_274_5267 <= 32'd0;
            operation_274_5266 <= 32'd0;
            operation_274_5265 <= 32'd0;
            operation_274_5264 <= 32'd0;
            operation_274_5263 <= 32'd0;
            operation_274_5262 <= 32'd0;
            operation_274_5261 <= 32'd0;
            operation_274_5260 <= 32'd0;
            operation_274_5259 <= 32'd0;
            operation_274_5258 <= 32'd0;
            operation_274_5257 <= 32'd0;
            operation_274_5332 <= 32'd0;
            operation_274_5331 <= 32'd0;
            operation_274_5330 <= 32'd0;
            operation_274_5329 <= 32'd0;
            operation_274_5328 <= 32'd0;
            operation_274_5327 <= 32'd0;
            operation_274_5326 <= 32'd0;
            operation_274_5325 <= 32'd0;
            operation_274_5324 <= 32'd0;
            operation_274_5323 <= 32'd0;
            operation_274_5322 <= 32'd0;
            operation_274_5321 <= 32'd0;
            operation_274_5320 <= 32'd0;
            operation_274_5319 <= 32'd0;
            operation_274_5318 <= 32'd0;
            operation_274_5317 <= 32'd0;
            operation_274_5352 <= 32'd0;
            operation_274_5351 <= 32'd0;
            operation_274_5350 <= 32'd0;
            operation_274_5349 <= 32'd0;
            operation_274_5348 <= 32'd0;
            operation_274_5347 <= 32'd0;
            operation_274_5346 <= 32'd0;
            operation_274_5345 <= 32'd0;
            operation_274_5344 <= 32'd0;
            operation_274_5343 <= 32'd0;
            operation_274_5342 <= 32'd0;
            operation_274_5341 <= 32'd0;
            operation_274_5340 <= 32'd0;
            operation_274_5339 <= 32'd0;
            operation_274_5338 <= 32'd0;
            operation_274_5337 <= 32'd0;
            operation_274_5376 <= 32'd0;
            operation_274_5375 <= 32'd0;
            operation_274_5374 <= 32'd0;
            operation_274_5373 <= 32'd0;
            operation_274_5372 <= 32'd0;
            operation_274_5371 <= 32'd0;
            operation_274_5370 <= 32'd0;
            operation_274_5369 <= 32'd0;
            operation_274_5368 <= 32'd0;
            operation_274_5367 <= 32'd0;
            operation_274_5366 <= 32'd0;
            operation_274_5365 <= 32'd0;
            operation_274_5364 <= 32'd0;
            operation_274_5363 <= 32'd0;
            operation_274_5362 <= 32'd0;
            operation_274_5361 <= 32'd0;
            operation_274_5414 <= 32'd0;
            operation_274_5413 <= 32'd0;
            operation_274_5412 <= 32'd0;
            operation_274_5411 <= 32'd0;
            operation_274_5410 <= 32'd0;
            operation_274_5409 <= 32'd0;
            operation_274_5408 <= 32'd0;
            operation_274_5407 <= 32'd0;
            operation_274_5406 <= 32'd0;
            operation_274_5405 <= 32'd0;
            operation_274_5404 <= 32'd0;
            operation_274_5403 <= 32'd0;
            operation_274_5402 <= 32'd0;
            operation_274_5401 <= 32'd0;
            operation_274_5400 <= 32'd0;
            operation_274_5399 <= 32'd0;
            operation_274_5398 <= 32'd0;
            operation_274_5397 <= 32'd0;
            operation_274_5396 <= 32'd0;
            operation_274_5395 <= 32'd0;
            operation_274_5394 <= 32'd0;
            operation_274_5393 <= 32'd0;
            operation_274_5392 <= 32'd0;
            operation_274_5391 <= 32'd0;
            operation_274_5390 <= 32'd0;
            operation_274_5389 <= 32'd0;
            operation_274_5388 <= 32'd0;
            operation_274_5387 <= 32'd0;
            operation_274_5386 <= 32'd0;
            operation_274_5385 <= 32'd0;
            operation_274_5384 <= 32'd0;
            operation_274_5383 <= 32'd0;
            operation_274_5440 <= 32'd0;
            operation_274_5439 <= 32'd0;
            operation_274_5422 <= 32'd0;
            operation_274_5421 <= 32'd0;
            operation_274_5464 <= 32'd0;
            operation_274_5463 <= 32'd0;
            operation_274_5446 <= 32'd0;
            operation_274_5445 <= 32'd0;
            operation_274_5485 <= 32'd0;
            operation_274_5484 <= 32'd0;
            operation_274_5483 <= 32'd0;
            operation_274_5482 <= 32'd0;
            operation_274_5481 <= 32'd0;
            operation_274_5480 <= 32'd0;
            operation_274_5479 <= 32'd0;
            operation_274_5478 <= 32'd0;
            operation_274_5477 <= 32'd0;
            operation_274_5476 <= 32'd0;
            operation_274_5475 <= 32'd0;
            operation_274_5474 <= 32'd0;
            operation_274_5473 <= 32'd0;
            operation_274_5472 <= 32'd0;
            operation_274_5471 <= 32'd0;
            operation_274_5470 <= 32'd0;
            operation_274_5536_latch <= 8'd0;
            operation_274_5535_latch <= 8'd0;
            operation_274_5534_latch <= 8'd0;
            operation_274_5533_latch <= 8'd0;
            operation_274_5532_latch <= 8'd0;
            operation_274_5531_latch <= 8'd0;
            operation_274_5530_latch <= 8'd0;
            operation_274_5529_latch <= 8'd0;
            operation_274_5528_latch <= 8'd0;
            operation_274_5527_latch <= 8'd0;
            operation_274_5526_latch <= 8'd0;
            operation_274_5525_latch <= 8'd0;
            operation_274_5524_latch <= 8'd0;
            operation_274_5523_latch <= 8'd0;
            operation_274_5522_latch <= 8'd0;
            operation_274_5521_latch <= 8'd0;
            operation_274_4733 <= 32'd0;
            operation_274_4732 <= 32'd0;
            operation_274_4731 <= 32'd0;
            operation_274_4730 <= 32'd0;
            operation_274_4729 <= 32'd0;
            operation_274_4728 <= 32'd0;
            operation_274_4727 <= 32'd0;
            operation_274_4726 <= 32'd0;
            operation_274_4725 <= 32'd0;
            operation_274_4724 <= 32'd0;
            operation_274_4723 <= 32'd0;
            operation_274_4722 <= 32'd0;
            operation_274_4721 <= 32'd0;
            operation_274_4720 <= 32'd0;
            operation_274_4719 <= 32'd0;
            operation_274_4718 <= 32'd0;
            operation_274_4785 <= 32'd0;
            operation_274_4784 <= 32'd0;
            operation_274_4783 <= 32'd0;
            operation_274_4782 <= 32'd0;
            operation_274_4781 <= 32'd0;
            operation_274_4780 <= 32'd0;
            operation_274_4779 <= 32'd0;
            operation_274_4778 <= 32'd0;
            operation_274_4777 <= 32'd0;
            operation_274_4776 <= 32'd0;
            operation_274_4775 <= 32'd0;
            operation_274_4774 <= 32'd0;
            operation_274_4773 <= 32'd0;
            operation_274_4772 <= 32'd0;
            operation_274_4771 <= 32'd0;
            operation_274_4770 <= 32'd0;
            operation_274_4843 <= 32'd0;
            operation_274_4842 <= 32'd0;
            operation_274_4841 <= 32'd0;
            operation_274_4840 <= 32'd0;
            operation_274_4839 <= 32'd0;
            operation_274_4838 <= 32'd0;
            operation_274_4837 <= 32'd0;
            operation_274_4836 <= 32'd0;
            operation_274_4835 <= 32'd0;
            operation_274_4834 <= 32'd0;
            operation_274_4833 <= 32'd0;
            operation_274_4832 <= 32'd0;
            operation_274_4831 <= 32'd0;
            operation_274_4830 <= 32'd0;
            operation_274_4829 <= 32'd0;
            operation_274_4828 <= 32'd0;
            operation_274_4903 <= 32'd0;
            operation_274_4902 <= 32'd0;
            operation_274_4901 <= 32'd0;
            operation_274_4900 <= 32'd0;
            operation_274_4899 <= 32'd0;
            operation_274_4898 <= 32'd0;
            operation_274_4897 <= 32'd0;
            operation_274_4896 <= 32'd0;
            operation_274_4895 <= 32'd0;
            operation_274_4894 <= 32'd0;
            operation_274_4893 <= 32'd0;
            operation_274_4892 <= 32'd0;
            operation_274_4891 <= 32'd0;
            operation_274_4890 <= 32'd0;
            operation_274_4889 <= 32'd0;
            operation_274_4888 <= 32'd0;
            operation_274_4923 <= 32'd0;
            operation_274_4922 <= 32'd0;
            operation_274_4921 <= 32'd0;
            operation_274_4920 <= 32'd0;
            operation_274_4919 <= 32'd0;
            operation_274_4918 <= 32'd0;
            operation_274_4917 <= 32'd0;
            operation_274_4916 <= 32'd0;
            operation_274_4915 <= 32'd0;
            operation_274_4914 <= 32'd0;
            operation_274_4913 <= 32'd0;
            operation_274_4912 <= 32'd0;
            operation_274_4911 <= 32'd0;
            operation_274_4910 <= 32'd0;
            operation_274_4909 <= 32'd0;
            operation_274_4908 <= 32'd0;
            operation_274_4947 <= 32'd0;
            operation_274_4946 <= 32'd0;
            operation_274_4945 <= 32'd0;
            operation_274_4944 <= 32'd0;
            operation_274_4943 <= 32'd0;
            operation_274_4942 <= 32'd0;
            operation_274_4941 <= 32'd0;
            operation_274_4940 <= 32'd0;
            operation_274_4939 <= 32'd0;
            operation_274_4938 <= 32'd0;
            operation_274_4937 <= 32'd0;
            operation_274_4936 <= 32'd0;
            operation_274_4935 <= 32'd0;
            operation_274_4934 <= 32'd0;
            operation_274_4933 <= 32'd0;
            operation_274_4932 <= 32'd0;
            operation_274_4985 <= 32'd0;
            operation_274_4984 <= 32'd0;
            operation_274_4983 <= 32'd0;
            operation_274_4982 <= 32'd0;
            operation_274_4981 <= 32'd0;
            operation_274_4980 <= 32'd0;
            operation_274_4979 <= 32'd0;
            operation_274_4978 <= 32'd0;
            operation_274_4977 <= 32'd0;
            operation_274_4976 <= 32'd0;
            operation_274_4975 <= 32'd0;
            operation_274_4974 <= 32'd0;
            operation_274_4973 <= 32'd0;
            operation_274_4972 <= 32'd0;
            operation_274_4971 <= 32'd0;
            operation_274_4970 <= 32'd0;
            operation_274_4969 <= 32'd0;
            operation_274_4968 <= 32'd0;
            operation_274_4967 <= 32'd0;
            operation_274_4966 <= 32'd0;
            operation_274_4965 <= 32'd0;
            operation_274_4964 <= 32'd0;
            operation_274_4963 <= 32'd0;
            operation_274_4962 <= 32'd0;
            operation_274_4961 <= 32'd0;
            operation_274_4960 <= 32'd0;
            operation_274_4959 <= 32'd0;
            operation_274_4958 <= 32'd0;
            operation_274_4957 <= 32'd0;
            operation_274_4956 <= 32'd0;
            operation_274_4955 <= 32'd0;
            operation_274_4954 <= 32'd0;
            operation_274_5011 <= 32'd0;
            operation_274_5010 <= 32'd0;
            operation_274_4993 <= 32'd0;
            operation_274_4992 <= 32'd0;
            operation_274_5035 <= 32'd0;
            operation_274_5034 <= 32'd0;
            operation_274_5017 <= 32'd0;
            operation_274_5016 <= 32'd0;
            operation_274_5056 <= 32'd0;
            operation_274_5055 <= 32'd0;
            operation_274_5054 <= 32'd0;
            operation_274_5053 <= 32'd0;
            operation_274_5052 <= 32'd0;
            operation_274_5051 <= 32'd0;
            operation_274_5050 <= 32'd0;
            operation_274_5049 <= 32'd0;
            operation_274_5048 <= 32'd0;
            operation_274_5047 <= 32'd0;
            operation_274_5046 <= 32'd0;
            operation_274_5045 <= 32'd0;
            operation_274_5044 <= 32'd0;
            operation_274_5043 <= 32'd0;
            operation_274_5042 <= 32'd0;
            operation_274_5041 <= 32'd0;
            operation_274_1536 <= 32'd0;
            operation_274_1560 <= 32'd0;
            operation_274_5107_latch <= 8'd0;
            operation_274_5106_latch <= 8'd0;
            operation_274_5105_latch <= 8'd0;
            operation_274_5104_latch <= 8'd0;
            operation_274_5103_latch <= 8'd0;
            operation_274_5102_latch <= 8'd0;
            operation_274_5101_latch <= 8'd0;
            operation_274_5100_latch <= 8'd0;
            operation_274_5099_latch <= 8'd0;
            operation_274_5098_latch <= 8'd0;
            operation_274_5097_latch <= 8'd0;
            operation_274_5096_latch <= 8'd0;
            operation_274_5095_latch <= 8'd0;
            operation_274_5094_latch <= 8'd0;
            operation_274_5093_latch <= 8'd0;
            operation_274_5092_latch <= 8'd0;
            operation_274_4304 <= 32'd0;
            operation_274_4303 <= 32'd0;
            operation_274_4302 <= 32'd0;
            operation_274_4301 <= 32'd0;
            operation_274_4300 <= 32'd0;
            operation_274_4299 <= 32'd0;
            operation_274_4298 <= 32'd0;
            operation_274_4297 <= 32'd0;
            operation_274_4296 <= 32'd0;
            operation_274_4295 <= 32'd0;
            operation_274_4294 <= 32'd0;
            operation_274_4293 <= 32'd0;
            operation_274_4292 <= 32'd0;
            operation_274_4291 <= 32'd0;
            operation_274_4290 <= 32'd0;
            operation_274_4289 <= 32'd0;
            operation_274_1544 <= 32'd0;
            operation_274_1504 <= 32'd0;
            operation_274_1552 <= 32'd0;
            operation_274_1528 <= 32'd0;
            operation_274_4356 <= 32'd0;
            operation_274_4355 <= 32'd0;
            operation_274_4354 <= 32'd0;
            operation_274_4353 <= 32'd0;
            operation_274_4352 <= 32'd0;
            operation_274_4351 <= 32'd0;
            operation_274_4350 <= 32'd0;
            operation_274_4349 <= 32'd0;
            operation_274_4348 <= 32'd0;
            operation_274_4347 <= 32'd0;
            operation_274_4346 <= 32'd0;
            operation_274_4345 <= 32'd0;
            operation_274_4344 <= 32'd0;
            operation_274_4343 <= 32'd0;
            operation_274_4342 <= 32'd0;
            operation_274_4341 <= 32'd0;
            operation_274_1512 <= 32'd0;
            operation_274_1472 <= 32'd0;
            operation_274_1520 <= 32'd0;
            operation_274_1496 <= 32'd0;
            operation_274_4414 <= 32'd0;
            operation_274_4413 <= 32'd0;
            operation_274_4412 <= 32'd0;
            operation_274_4411 <= 32'd0;
            operation_274_4410 <= 32'd0;
            operation_274_4409 <= 32'd0;
            operation_274_4408 <= 32'd0;
            operation_274_4407 <= 32'd0;
            operation_274_4406 <= 32'd0;
            operation_274_4405 <= 32'd0;
            operation_274_4404 <= 32'd0;
            operation_274_4403 <= 32'd0;
            operation_274_4402 <= 32'd0;
            operation_274_4401 <= 32'd0;
            operation_274_4400 <= 32'd0;
            operation_274_4399 <= 32'd0;
            operation_274_1480 <= 32'd0;
            operation_274_1440 <= 32'd0;
            operation_274_1488 <= 32'd0;
            operation_274_1464 <= 32'd0;
            operation_274_1423_latch <= 8'd0;
            operation_274_4474 <= 32'd0;
            operation_274_4473 <= 32'd0;
            operation_274_4472 <= 32'd0;
            operation_274_4471 <= 32'd0;
            operation_274_4470 <= 32'd0;
            operation_274_4469 <= 32'd0;
            operation_274_4468 <= 32'd0;
            operation_274_4467 <= 32'd0;
            operation_274_4466 <= 32'd0;
            operation_274_4465 <= 32'd0;
            operation_274_4464 <= 32'd0;
            operation_274_4463 <= 32'd0;
            operation_274_4462 <= 32'd0;
            operation_274_4461 <= 32'd0;
            operation_274_4460 <= 32'd0;
            operation_274_4459 <= 32'd0;
            operation_274_1448 <= 32'd0;
            operation_274_1432 <= 32'd0;
            operation_274_1456 <= 32'd0;
            operation_274_4494 <= 32'd0;
            operation_274_4493 <= 32'd0;
            operation_274_4492 <= 32'd0;
            operation_274_4491 <= 32'd0;
            operation_274_4490 <= 32'd0;
            operation_274_4489 <= 32'd0;
            operation_274_4488 <= 32'd0;
            operation_274_4487 <= 32'd0;
            operation_274_4486 <= 32'd0;
            operation_274_4485 <= 32'd0;
            operation_274_4484 <= 32'd0;
            operation_274_4483 <= 32'd0;
            operation_274_4482 <= 32'd0;
            operation_274_4481 <= 32'd0;
            operation_274_4480 <= 32'd0;
            operation_274_4479 <= 32'd0;
            operation_274_5198 <= 32'd0;
            operation_274_4518 <= 32'd0;
            operation_274_4517 <= 32'd0;
            operation_274_4516 <= 32'd0;
            operation_274_4515 <= 32'd0;
            operation_274_4514 <= 32'd0;
            operation_274_4513 <= 32'd0;
            operation_274_4512 <= 32'd0;
            operation_274_4511 <= 32'd0;
            operation_274_4510 <= 32'd0;
            operation_274_4509 <= 32'd0;
            operation_274_4508 <= 32'd0;
            operation_274_4507 <= 32'd0;
            operation_274_4506 <= 32'd0;
            operation_274_4505 <= 32'd0;
            operation_274_4504 <= 32'd0;
            operation_274_4503 <= 32'd0;
            operation_274_1418_latch <= 8'd0;
            operation_274_1408_latch <= 8'd0;
            operation_274_1413_latch <= 8'd0;
            operation_274_4556 <= 32'd0;
            operation_274_4555 <= 32'd0;
            operation_274_4554 <= 32'd0;
            operation_274_4553 <= 32'd0;
            operation_274_4552 <= 32'd0;
            operation_274_4551 <= 32'd0;
            operation_274_4550 <= 32'd0;
            operation_274_4549 <= 32'd0;
            operation_274_4548 <= 32'd0;
            operation_274_4547 <= 32'd0;
            operation_274_4546 <= 32'd0;
            operation_274_4545 <= 32'd0;
            operation_274_4544 <= 32'd0;
            operation_274_4543 <= 32'd0;
            operation_274_4542 <= 32'd0;
            operation_274_4541 <= 32'd0;
            operation_274_4540 <= 32'd0;
            operation_274_4539 <= 32'd0;
            operation_274_4538 <= 32'd0;
            operation_274_4537 <= 32'd0;
            operation_274_4536 <= 32'd0;
            operation_274_4535 <= 32'd0;
            operation_274_4534 <= 32'd0;
            operation_274_4533 <= 32'd0;
            operation_274_4532 <= 32'd0;
            operation_274_4531 <= 32'd0;
            operation_274_4530 <= 32'd0;
            operation_274_4529 <= 32'd0;
            operation_274_4528 <= 32'd0;
            operation_274_4527 <= 32'd0;
            operation_274_4526 <= 32'd0;
            operation_274_4525 <= 32'd0;
            operation_274_4582 <= 32'd0;
            operation_274_4581 <= 32'd0;
            operation_274_4564 <= 32'd0;
            operation_274_4563 <= 32'd0;
            operation_274_5274 <= 32'd0;
            operation_274_5273 <= 32'd0;
            operation_274_5256 <= 32'd0;
            operation_274_5255 <= 32'd0;
            operation_274_4606 <= 32'd0;
            operation_274_4605 <= 32'd0;
            operation_274_4588 <= 32'd0;
            operation_274_4587 <= 32'd0;
            operation_274_4627 <= 32'd0;
            operation_274_4626 <= 32'd0;
            operation_274_4625 <= 32'd0;
            operation_274_4624 <= 32'd0;
            operation_274_4623 <= 32'd0;
            operation_274_4622 <= 32'd0;
            operation_274_4621 <= 32'd0;
            operation_274_4620 <= 32'd0;
            operation_274_4619 <= 32'd0;
            operation_274_4618 <= 32'd0;
            operation_274_4617 <= 32'd0;
            operation_274_4616 <= 32'd0;
            operation_274_4615 <= 32'd0;
            operation_274_4614 <= 32'd0;
            operation_274_4613 <= 32'd0;
            operation_274_4612 <= 32'd0;
            operation_274_5334 <= 32'd0;
            operation_274_5333 <= 32'd0;
            operation_274_5316 <= 32'd0;
            operation_274_5315 <= 32'd0;
            operation_274_4678_latch <= 8'd0;
            operation_274_4677_latch <= 8'd0;
            operation_274_4676_latch <= 8'd0;
            operation_274_4675_latch <= 8'd0;
            operation_274_4674_latch <= 8'd0;
            operation_274_4673_latch <= 8'd0;
            operation_274_4672_latch <= 8'd0;
            operation_274_4671_latch <= 8'd0;
            operation_274_4670_latch <= 8'd0;
            operation_274_4669_latch <= 8'd0;
            operation_274_4668_latch <= 8'd0;
            operation_274_4667_latch <= 8'd0;
            operation_274_4666_latch <= 8'd0;
            operation_274_4665_latch <= 8'd0;
            operation_274_4664_latch <= 8'd0;
            operation_274_4663_latch <= 8'd0;
            operation_274_3875 <= 32'd0;
            operation_274_3874 <= 32'd0;
            operation_274_3873 <= 32'd0;
            operation_274_3872 <= 32'd0;
            operation_274_3871 <= 32'd0;
            operation_274_3870 <= 32'd0;
            operation_274_3869 <= 32'd0;
            operation_274_3868 <= 32'd0;
            operation_274_3867 <= 32'd0;
            operation_274_3866 <= 32'd0;
            operation_274_3865 <= 32'd0;
            operation_274_3864 <= 32'd0;
            operation_274_3863 <= 32'd0;
            operation_274_3862 <= 32'd0;
            operation_274_3861 <= 32'd0;
            operation_274_3860 <= 32'd0;
            operation_274_5418 <= 32'd0;
            operation_274_5417 <= 32'd0;
            operation_274_5380 <= 32'd0;
            operation_274_5379 <= 32'd0;
            operation_274_3927 <= 32'd0;
            operation_274_3926 <= 32'd0;
            operation_274_3925 <= 32'd0;
            operation_274_3924 <= 32'd0;
            operation_274_3923 <= 32'd0;
            operation_274_3922 <= 32'd0;
            operation_274_3921 <= 32'd0;
            operation_274_3920 <= 32'd0;
            operation_274_3919 <= 32'd0;
            operation_274_3918 <= 32'd0;
            operation_274_3917 <= 32'd0;
            operation_274_3916 <= 32'd0;
            operation_274_3915 <= 32'd0;
            operation_274_3914 <= 32'd0;
            operation_274_3913 <= 32'd0;
            operation_274_3912 <= 32'd0;
            operation_274_5488 <= 32'd0;
            operation_274_5487 <= 32'd0;
            operation_274_5486 <= 32'd0;
            operation_274_5469 <= 32'd0;
            operation_274_5538_latch <= 8'd0;
            operation_274_5537_latch <= 8'd0;
            operation_274_5520_latch <= 8'd0;
            operation_274_5519_latch <= 8'd0;
            operation_274_3985 <= 32'd0;
            operation_274_3984 <= 32'd0;
            operation_274_3983 <= 32'd0;
            operation_274_3982 <= 32'd0;
            operation_274_3981 <= 32'd0;
            operation_274_3980 <= 32'd0;
            operation_274_3979 <= 32'd0;
            operation_274_3978 <= 32'd0;
            operation_274_3977 <= 32'd0;
            operation_274_3976 <= 32'd0;
            operation_274_3975 <= 32'd0;
            operation_274_3974 <= 32'd0;
            operation_274_3973 <= 32'd0;
            operation_274_3972 <= 32'd0;
            operation_274_3971 <= 32'd0;
            operation_274_3970 <= 32'd0;
            operation_274_4845 <= 32'd0;
            operation_274_4844 <= 32'd0;
            operation_274_4826 <= 32'd0;
            operation_274_4769 <= 32'd0;
            operation_274_4045 <= 32'd0;
            operation_274_4044 <= 32'd0;
            operation_274_4043 <= 32'd0;
            operation_274_4042 <= 32'd0;
            operation_274_4041 <= 32'd0;
            operation_274_4040 <= 32'd0;
            operation_274_4039 <= 32'd0;
            operation_274_4038 <= 32'd0;
            operation_274_4037 <= 32'd0;
            operation_274_4036 <= 32'd0;
            operation_274_4035 <= 32'd0;
            operation_274_4034 <= 32'd0;
            operation_274_4033 <= 32'd0;
            operation_274_4032 <= 32'd0;
            operation_274_4031 <= 32'd0;
            operation_274_4030 <= 32'd0;
            operation_274_4065 <= 32'd0;
            operation_274_4064 <= 32'd0;
            operation_274_4063 <= 32'd0;
            operation_274_4062 <= 32'd0;
            operation_274_4061 <= 32'd0;
            operation_274_4060 <= 32'd0;
            operation_274_4059 <= 32'd0;
            operation_274_4058 <= 32'd0;
            operation_274_4057 <= 32'd0;
            operation_274_4056 <= 32'd0;
            operation_274_4055 <= 32'd0;
            operation_274_4054 <= 32'd0;
            operation_274_4053 <= 32'd0;
            operation_274_4052 <= 32'd0;
            operation_274_4051 <= 32'd0;
            operation_274_4050 <= 32'd0;
            operation_274_4905 <= 32'd0;
            operation_274_4904 <= 32'd0;
            operation_274_4886 <= 32'd0;
            operation_274_4827 <= 32'd0;
            operation_274_4089 <= 32'd0;
            operation_274_4088 <= 32'd0;
            operation_274_4087 <= 32'd0;
            operation_274_4086 <= 32'd0;
            operation_274_4085 <= 32'd0;
            operation_274_4084 <= 32'd0;
            operation_274_4083 <= 32'd0;
            operation_274_4082 <= 32'd0;
            operation_274_4081 <= 32'd0;
            operation_274_4080 <= 32'd0;
            operation_274_4079 <= 32'd0;
            operation_274_4078 <= 32'd0;
            operation_274_4077 <= 32'd0;
            operation_274_4076 <= 32'd0;
            operation_274_4075 <= 32'd0;
            operation_274_4074 <= 32'd0;
            operation_274_4127 <= 32'd0;
            operation_274_4126 <= 32'd0;
            operation_274_4125 <= 32'd0;
            operation_274_4124 <= 32'd0;
            operation_274_4123 <= 32'd0;
            operation_274_4122 <= 32'd0;
            operation_274_4121 <= 32'd0;
            operation_274_4120 <= 32'd0;
            operation_274_4119 <= 32'd0;
            operation_274_4118 <= 32'd0;
            operation_274_4117 <= 32'd0;
            operation_274_4116 <= 32'd0;
            operation_274_4115 <= 32'd0;
            operation_274_4114 <= 32'd0;
            operation_274_4113 <= 32'd0;
            operation_274_4112 <= 32'd0;
            operation_274_4111 <= 32'd0;
            operation_274_4110 <= 32'd0;
            operation_274_4109 <= 32'd0;
            operation_274_4108 <= 32'd0;
            operation_274_4107 <= 32'd0;
            operation_274_4106 <= 32'd0;
            operation_274_4105 <= 32'd0;
            operation_274_4104 <= 32'd0;
            operation_274_4103 <= 32'd0;
            operation_274_4102 <= 32'd0;
            operation_274_4101 <= 32'd0;
            operation_274_4100 <= 32'd0;
            operation_274_4099 <= 32'd0;
            operation_274_4098 <= 32'd0;
            operation_274_4097 <= 32'd0;
            operation_274_4096 <= 32'd0;
            operation_274_4153 <= 32'd0;
            operation_274_4152 <= 32'd0;
            operation_274_4135 <= 32'd0;
            operation_274_4134 <= 32'd0;
            operation_274_4989 <= 32'd0;
            operation_274_4988 <= 32'd0;
            operation_274_4950 <= 32'd0;
            operation_274_4887 <= 32'd0;
            operation_274_4177 <= 32'd0;
            operation_274_4176 <= 32'd0;
            operation_274_4159 <= 32'd0;
            operation_274_4158 <= 32'd0;
            operation_274_4198 <= 32'd0;
            operation_274_4197 <= 32'd0;
            operation_274_4196 <= 32'd0;
            operation_274_4195 <= 32'd0;
            operation_274_4194 <= 32'd0;
            operation_274_4193 <= 32'd0;
            operation_274_4192 <= 32'd0;
            operation_274_4191 <= 32'd0;
            operation_274_4190 <= 32'd0;
            operation_274_4189 <= 32'd0;
            operation_274_4188 <= 32'd0;
            operation_274_4187 <= 32'd0;
            operation_274_4186 <= 32'd0;
            operation_274_4185 <= 32'd0;
            operation_274_4184 <= 32'd0;
            operation_274_4183 <= 32'd0;
            operation_274_5059 <= 32'd0;
            operation_274_5058 <= 32'd0;
            operation_274_5040 <= 32'd0;
            operation_274_4951 <= 32'd0;
            operation_274_4249_latch <= 8'd0;
            operation_274_4248_latch <= 8'd0;
            operation_274_4247_latch <= 8'd0;
            operation_274_4246_latch <= 8'd0;
            operation_274_4245_latch <= 8'd0;
            operation_274_4244_latch <= 8'd0;
            operation_274_4243_latch <= 8'd0;
            operation_274_4242_latch <= 8'd0;
            operation_274_4241_latch <= 8'd0;
            operation_274_4240_latch <= 8'd0;
            operation_274_4239_latch <= 8'd0;
            operation_274_4238_latch <= 8'd0;
            operation_274_4237_latch <= 8'd0;
            operation_274_4236_latch <= 8'd0;
            operation_274_4235_latch <= 8'd0;
            operation_274_4234_latch <= 8'd0;
            operation_274_5109_latch <= 8'd0;
            operation_274_5091_latch <= 8'd0;
            operation_274_5090_latch <= 8'd0;
            operation_274_3446 <= 32'd0;
            operation_274_3445 <= 32'd0;
            operation_274_3444 <= 32'd0;
            operation_274_3443 <= 32'd0;
            operation_274_3442 <= 32'd0;
            operation_274_3441 <= 32'd0;
            operation_274_3440 <= 32'd0;
            operation_274_3439 <= 32'd0;
            operation_274_3438 <= 32'd0;
            operation_274_3437 <= 32'd0;
            operation_274_3436 <= 32'd0;
            operation_274_3435 <= 32'd0;
            operation_274_3434 <= 32'd0;
            operation_274_3433 <= 32'd0;
            operation_274_3432 <= 32'd0;
            operation_274_3431 <= 32'd0;
            operation_274_5057 <= 32'd0;
            operation_274_4416 <= 32'd0;
            operation_274_4397 <= 32'd0;
            operation_274_4340 <= 32'd0;
            operation_274_5108_latch <= 8'd0;
            operation_274_3498 <= 32'd0;
            operation_274_3497 <= 32'd0;
            operation_274_3496 <= 32'd0;
            operation_274_3495 <= 32'd0;
            operation_274_3494 <= 32'd0;
            operation_274_3493 <= 32'd0;
            operation_274_3492 <= 32'd0;
            operation_274_3491 <= 32'd0;
            operation_274_3490 <= 32'd0;
            operation_274_3489 <= 32'd0;
            operation_274_3488 <= 32'd0;
            operation_274_3487 <= 32'd0;
            operation_274_3486 <= 32'd0;
            operation_274_3485 <= 32'd0;
            operation_274_3484 <= 32'd0;
            operation_274_3483 <= 32'd0;
            operation_274_4476 <= 32'd0;
            operation_274_4457 <= 32'd0;
            operation_274_4415 <= 32'd0;
            operation_274_4398 <= 32'd0;
            operation_274_3556 <= 32'd0;
            operation_274_3555 <= 32'd0;
            operation_274_3554 <= 32'd0;
            operation_274_3553 <= 32'd0;
            operation_274_3552 <= 32'd0;
            operation_274_3551 <= 32'd0;
            operation_274_3550 <= 32'd0;
            operation_274_3549 <= 32'd0;
            operation_274_3548 <= 32'd0;
            operation_274_3547 <= 32'd0;
            operation_274_3546 <= 32'd0;
            operation_274_3545 <= 32'd0;
            operation_274_3544 <= 32'd0;
            operation_274_3543 <= 32'd0;
            operation_274_3542 <= 32'd0;
            operation_274_3541 <= 32'd0;
            operation_274_4560 <= 32'd0;
            operation_274_4521 <= 32'd0;
            operation_274_4475 <= 32'd0;
            operation_274_4458 <= 32'd0;
            operation_274_3616 <= 32'd0;
            operation_274_3615 <= 32'd0;
            operation_274_3614 <= 32'd0;
            operation_274_3613 <= 32'd0;
            operation_274_3612 <= 32'd0;
            operation_274_3611 <= 32'd0;
            operation_274_3610 <= 32'd0;
            operation_274_3609 <= 32'd0;
            operation_274_3608 <= 32'd0;
            operation_274_3607 <= 32'd0;
            operation_274_3606 <= 32'd0;
            operation_274_3605 <= 32'd0;
            operation_274_3604 <= 32'd0;
            operation_274_3603 <= 32'd0;
            operation_274_3602 <= 32'd0;
            operation_274_3601 <= 32'd0;
            operation_274_3636 <= 32'd0;
            operation_274_3635 <= 32'd0;
            operation_274_3634 <= 32'd0;
            operation_274_3633 <= 32'd0;
            operation_274_3632 <= 32'd0;
            operation_274_3631 <= 32'd0;
            operation_274_3630 <= 32'd0;
            operation_274_3629 <= 32'd0;
            operation_274_3628 <= 32'd0;
            operation_274_3627 <= 32'd0;
            operation_274_3626 <= 32'd0;
            operation_274_3625 <= 32'd0;
            operation_274_3624 <= 32'd0;
            operation_274_3623 <= 32'd0;
            operation_274_3622 <= 32'd0;
            operation_274_3621 <= 32'd0;
            operation_274_4630 <= 32'd0;
            operation_274_4611 <= 32'd0;
            operation_274_4559 <= 32'd0;
            operation_274_4522 <= 32'd0;
            operation_274_3660 <= 32'd0;
            operation_274_3659 <= 32'd0;
            operation_274_3658 <= 32'd0;
            operation_274_3657 <= 32'd0;
            operation_274_3656 <= 32'd0;
            operation_274_3655 <= 32'd0;
            operation_274_3654 <= 32'd0;
            operation_274_3653 <= 32'd0;
            operation_274_3652 <= 32'd0;
            operation_274_3651 <= 32'd0;
            operation_274_3650 <= 32'd0;
            operation_274_3649 <= 32'd0;
            operation_274_3648 <= 32'd0;
            operation_274_3647 <= 32'd0;
            operation_274_3646 <= 32'd0;
            operation_274_3645 <= 32'd0;
            operation_274_3698 <= 32'd0;
            operation_274_3697 <= 32'd0;
            operation_274_3696 <= 32'd0;
            operation_274_3695 <= 32'd0;
            operation_274_3694 <= 32'd0;
            operation_274_3693 <= 32'd0;
            operation_274_3692 <= 32'd0;
            operation_274_3691 <= 32'd0;
            operation_274_3690 <= 32'd0;
            operation_274_3689 <= 32'd0;
            operation_274_3688 <= 32'd0;
            operation_274_3687 <= 32'd0;
            operation_274_3686 <= 32'd0;
            operation_274_3685 <= 32'd0;
            operation_274_3684 <= 32'd0;
            operation_274_3683 <= 32'd0;
            operation_274_3682 <= 32'd0;
            operation_274_3681 <= 32'd0;
            operation_274_3680 <= 32'd0;
            operation_274_3679 <= 32'd0;
            operation_274_3678 <= 32'd0;
            operation_274_3677 <= 32'd0;
            operation_274_3676 <= 32'd0;
            operation_274_3675 <= 32'd0;
            operation_274_3674 <= 32'd0;
            operation_274_3673 <= 32'd0;
            operation_274_3672 <= 32'd0;
            operation_274_3671 <= 32'd0;
            operation_274_3670 <= 32'd0;
            operation_274_3669 <= 32'd0;
            operation_274_3668 <= 32'd0;
            operation_274_3667 <= 32'd0;
            operation_274_4680_latch <= 8'd0;
            operation_274_4661_latch <= 8'd0;
            operation_274_3724 <= 32'd0;
            operation_274_3723 <= 32'd0;
            operation_274_3706 <= 32'd0;
            operation_274_3705 <= 32'd0;
            operation_274_4629 <= 32'd0;
            operation_274_4628 <= 32'd0;
            operation_274_3748 <= 32'd0;
            operation_274_3747 <= 32'd0;
            operation_274_3730 <= 32'd0;
            operation_274_3729 <= 32'd0;
            operation_274_3987 <= 32'd0;
            operation_274_3911 <= 32'd0;
            operation_274_3769 <= 32'd0;
            operation_274_3768 <= 32'd0;
            operation_274_3767 <= 32'd0;
            operation_274_3766 <= 32'd0;
            operation_274_3765 <= 32'd0;
            operation_274_3764 <= 32'd0;
            operation_274_3763 <= 32'd0;
            operation_274_3762 <= 32'd0;
            operation_274_3761 <= 32'd0;
            operation_274_3760 <= 32'd0;
            operation_274_3759 <= 32'd0;
            operation_274_3758 <= 32'd0;
            operation_274_3757 <= 32'd0;
            operation_274_3756 <= 32'd0;
            operation_274_3755 <= 32'd0;
            operation_274_3754 <= 32'd0;
            operation_274_4679_latch <= 8'd0;
            operation_274_4662_latch <= 8'd0;
            operation_274_3820_latch <= 8'd0;
            operation_274_3819_latch <= 8'd0;
            operation_274_3818_latch <= 8'd0;
            operation_274_3817_latch <= 8'd0;
            operation_274_3816_latch <= 8'd0;
            operation_274_3815_latch <= 8'd0;
            operation_274_3814_latch <= 8'd0;
            operation_274_3813_latch <= 8'd0;
            operation_274_3812_latch <= 8'd0;
            operation_274_3811_latch <= 8'd0;
            operation_274_3810_latch <= 8'd0;
            operation_274_3809_latch <= 8'd0;
            operation_274_3808_latch <= 8'd0;
            operation_274_3807_latch <= 8'd0;
            operation_274_3806_latch <= 8'd0;
            operation_274_3805_latch <= 8'd0;
            operation_274_4047 <= 32'd0;
            operation_274_3986 <= 32'd0;
            operation_274_3969 <= 32'd0;
            operation_274_3968 <= 32'd0;
            operation_274_3017 <= 32'd0;
            operation_274_3016 <= 32'd0;
            operation_274_3015 <= 32'd0;
            operation_274_3014 <= 32'd0;
            operation_274_3013 <= 32'd0;
            operation_274_3012 <= 32'd0;
            operation_274_3011 <= 32'd0;
            operation_274_3010 <= 32'd0;
            operation_274_3009 <= 32'd0;
            operation_274_3008 <= 32'd0;
            operation_274_3007 <= 32'd0;
            operation_274_3006 <= 32'd0;
            operation_274_3005 <= 32'd0;
            operation_274_3004 <= 32'd0;
            operation_274_3003 <= 32'd0;
            operation_274_3002 <= 32'd0;
            operation_274_4131 <= 32'd0;
            operation_274_4046 <= 32'd0;
            operation_274_4029 <= 32'd0;
            operation_274_4028 <= 32'd0;
            operation_274_3069 <= 32'd0;
            operation_274_3068 <= 32'd0;
            operation_274_3067 <= 32'd0;
            operation_274_3066 <= 32'd0;
            operation_274_3065 <= 32'd0;
            operation_274_3064 <= 32'd0;
            operation_274_3063 <= 32'd0;
            operation_274_3062 <= 32'd0;
            operation_274_3061 <= 32'd0;
            operation_274_3060 <= 32'd0;
            operation_274_3059 <= 32'd0;
            operation_274_3058 <= 32'd0;
            operation_274_3057 <= 32'd0;
            operation_274_3056 <= 32'd0;
            operation_274_3055 <= 32'd0;
            operation_274_3054 <= 32'd0;
            operation_274_4201 <= 32'd0;
            operation_274_4130 <= 32'd0;
            operation_274_4093 <= 32'd0;
            operation_274_4092 <= 32'd0;
            operation_274_3127 <= 32'd0;
            operation_274_3126 <= 32'd0;
            operation_274_3125 <= 32'd0;
            operation_274_3124 <= 32'd0;
            operation_274_3123 <= 32'd0;
            operation_274_3122 <= 32'd0;
            operation_274_3121 <= 32'd0;
            operation_274_3120 <= 32'd0;
            operation_274_3119 <= 32'd0;
            operation_274_3118 <= 32'd0;
            operation_274_3117 <= 32'd0;
            operation_274_3116 <= 32'd0;
            operation_274_3115 <= 32'd0;
            operation_274_3114 <= 32'd0;
            operation_274_3113 <= 32'd0;
            operation_274_3112 <= 32'd0;
            operation_274_4232_latch <= 8'd0;
            operation_274_4200 <= 32'd0;
            operation_274_4199 <= 32'd0;
            operation_274_4182 <= 32'd0;
            operation_274_3482 <= 32'd0;
            operation_274_3187 <= 32'd0;
            operation_274_3186 <= 32'd0;
            operation_274_3185 <= 32'd0;
            operation_274_3184 <= 32'd0;
            operation_274_3183 <= 32'd0;
            operation_274_3182 <= 32'd0;
            operation_274_3181 <= 32'd0;
            operation_274_3180 <= 32'd0;
            operation_274_3179 <= 32'd0;
            operation_274_3178 <= 32'd0;
            operation_274_3177 <= 32'd0;
            operation_274_3176 <= 32'd0;
            operation_274_3175 <= 32'd0;
            operation_274_3174 <= 32'd0;
            operation_274_3173 <= 32'd0;
            operation_274_3172 <= 32'd0;
            operation_274_4251_latch <= 8'd0;
            operation_274_4250_latch <= 8'd0;
            operation_274_4233_latch <= 8'd0;
            operation_274_3207 <= 32'd0;
            operation_274_3206 <= 32'd0;
            operation_274_3205 <= 32'd0;
            operation_274_3204 <= 32'd0;
            operation_274_3203 <= 32'd0;
            operation_274_3202 <= 32'd0;
            operation_274_3201 <= 32'd0;
            operation_274_3200 <= 32'd0;
            operation_274_3199 <= 32'd0;
            operation_274_3198 <= 32'd0;
            operation_274_3197 <= 32'd0;
            operation_274_3196 <= 32'd0;
            operation_274_3195 <= 32'd0;
            operation_274_3194 <= 32'd0;
            operation_274_3193 <= 32'd0;
            operation_274_3192 <= 32'd0;
            operation_274_3231 <= 32'd0;
            operation_274_3230 <= 32'd0;
            operation_274_3229 <= 32'd0;
            operation_274_3228 <= 32'd0;
            operation_274_3227 <= 32'd0;
            operation_274_3226 <= 32'd0;
            operation_274_3225 <= 32'd0;
            operation_274_3224 <= 32'd0;
            operation_274_3223 <= 32'd0;
            operation_274_3222 <= 32'd0;
            operation_274_3221 <= 32'd0;
            operation_274_3220 <= 32'd0;
            operation_274_3219 <= 32'd0;
            operation_274_3218 <= 32'd0;
            operation_274_3217 <= 32'd0;
            operation_274_3216 <= 32'd0;
            operation_274_3558 <= 32'd0;
            operation_274_3557 <= 32'd0;
            operation_274_3540 <= 32'd0;
            operation_274_3539 <= 32'd0;
            operation_274_3269 <= 32'd0;
            operation_274_3268 <= 32'd0;
            operation_274_3267 <= 32'd0;
            operation_274_3266 <= 32'd0;
            operation_274_3265 <= 32'd0;
            operation_274_3264 <= 32'd0;
            operation_274_3263 <= 32'd0;
            operation_274_3262 <= 32'd0;
            operation_274_3261 <= 32'd0;
            operation_274_3260 <= 32'd0;
            operation_274_3259 <= 32'd0;
            operation_274_3258 <= 32'd0;
            operation_274_3257 <= 32'd0;
            operation_274_3256 <= 32'd0;
            operation_274_3255 <= 32'd0;
            operation_274_3254 <= 32'd0;
            operation_274_3253 <= 32'd0;
            operation_274_3252 <= 32'd0;
            operation_274_3251 <= 32'd0;
            operation_274_3250 <= 32'd0;
            operation_274_3249 <= 32'd0;
            operation_274_3248 <= 32'd0;
            operation_274_3247 <= 32'd0;
            operation_274_3246 <= 32'd0;
            operation_274_3245 <= 32'd0;
            operation_274_3244 <= 32'd0;
            operation_274_3243 <= 32'd0;
            operation_274_3242 <= 32'd0;
            operation_274_3241 <= 32'd0;
            operation_274_3240 <= 32'd0;
            operation_274_3239 <= 32'd0;
            operation_274_3238 <= 32'd0;
            operation_274_3295 <= 32'd0;
            operation_274_3294 <= 32'd0;
            operation_274_3277 <= 32'd0;
            operation_274_3276 <= 32'd0;
            operation_274_3319 <= 32'd0;
            operation_274_3318 <= 32'd0;
            operation_274_3301 <= 32'd0;
            operation_274_3300 <= 32'd0;
            operation_274_3618 <= 32'd0;
            operation_274_3617 <= 32'd0;
            operation_274_3600 <= 32'd0;
            operation_274_3599 <= 32'd0;
            operation_274_3340 <= 32'd0;
            operation_274_3339 <= 32'd0;
            operation_274_3338 <= 32'd0;
            operation_274_3337 <= 32'd0;
            operation_274_3336 <= 32'd0;
            operation_274_3335 <= 32'd0;
            operation_274_3334 <= 32'd0;
            operation_274_3333 <= 32'd0;
            operation_274_3332 <= 32'd0;
            operation_274_3331 <= 32'd0;
            operation_274_3330 <= 32'd0;
            operation_274_3329 <= 32'd0;
            operation_274_3328 <= 32'd0;
            operation_274_3327 <= 32'd0;
            operation_274_3326 <= 32'd0;
            operation_274_3325 <= 32'd0;
            operation_274_3391_latch <= 8'd0;
            operation_274_3390_latch <= 8'd0;
            operation_274_3389_latch <= 8'd0;
            operation_274_3388_latch <= 8'd0;
            operation_274_3387_latch <= 8'd0;
            operation_274_3386_latch <= 8'd0;
            operation_274_3385_latch <= 8'd0;
            operation_274_3384_latch <= 8'd0;
            operation_274_3383_latch <= 8'd0;
            operation_274_3382_latch <= 8'd0;
            operation_274_3381_latch <= 8'd0;
            operation_274_3380_latch <= 8'd0;
            operation_274_3379_latch <= 8'd0;
            operation_274_3378_latch <= 8'd0;
            operation_274_3377_latch <= 8'd0;
            operation_274_3376_latch <= 8'd0;
            operation_274_3702 <= 32'd0;
            operation_274_3701 <= 32'd0;
            operation_274_3664 <= 32'd0;
            operation_274_3663 <= 32'd0;
            operation_274_2588 <= 32'd0;
            operation_274_2587 <= 32'd0;
            operation_274_2586 <= 32'd0;
            operation_274_2585 <= 32'd0;
            operation_274_2584 <= 32'd0;
            operation_274_2583 <= 32'd0;
            operation_274_2582 <= 32'd0;
            operation_274_2581 <= 32'd0;
            operation_274_2580 <= 32'd0;
            operation_274_2579 <= 32'd0;
            operation_274_2578 <= 32'd0;
            operation_274_2577 <= 32'd0;
            operation_274_2576 <= 32'd0;
            operation_274_2575 <= 32'd0;
            operation_274_2574 <= 32'd0;
            operation_274_2573 <= 32'd0;
            operation_274_3772 <= 32'd0;
            operation_274_3771 <= 32'd0;
            operation_274_3770 <= 32'd0;
            operation_274_3753 <= 32'd0;
            operation_274_2640 <= 32'd0;
            operation_274_2639 <= 32'd0;
            operation_274_2638 <= 32'd0;
            operation_274_2637 <= 32'd0;
            operation_274_2636 <= 32'd0;
            operation_274_2635 <= 32'd0;
            operation_274_2634 <= 32'd0;
            operation_274_2633 <= 32'd0;
            operation_274_2632 <= 32'd0;
            operation_274_2631 <= 32'd0;
            operation_274_2630 <= 32'd0;
            operation_274_2629 <= 32'd0;
            operation_274_2628 <= 32'd0;
            operation_274_2627 <= 32'd0;
            operation_274_2626 <= 32'd0;
            operation_274_2625 <= 32'd0;
            operation_274_3822_latch <= 8'd0;
            operation_274_3821_latch <= 8'd0;
            operation_274_3804_latch <= 8'd0;
            operation_274_3803_latch <= 8'd0;
            operation_274_3129 <= 32'd0;
            operation_274_3128 <= 32'd0;
            operation_274_3110 <= 32'd0;
            operation_274_3053 <= 32'd0;
            operation_274_2698 <= 32'd0;
            operation_274_2697 <= 32'd0;
            operation_274_2696 <= 32'd0;
            operation_274_2695 <= 32'd0;
            operation_274_2694 <= 32'd0;
            operation_274_2693 <= 32'd0;
            operation_274_2692 <= 32'd0;
            operation_274_2691 <= 32'd0;
            operation_274_2690 <= 32'd0;
            operation_274_2689 <= 32'd0;
            operation_274_2688 <= 32'd0;
            operation_274_2687 <= 32'd0;
            operation_274_2686 <= 32'd0;
            operation_274_2685 <= 32'd0;
            operation_274_2684 <= 32'd0;
            operation_274_2683 <= 32'd0;
            operation_274_3189 <= 32'd0;
            operation_274_3188 <= 32'd0;
            operation_274_3170 <= 32'd0;
            operation_274_3111 <= 32'd0;
            operation_274_2758 <= 32'd0;
            operation_274_2757 <= 32'd0;
            operation_274_2756 <= 32'd0;
            operation_274_2755 <= 32'd0;
            operation_274_2754 <= 32'd0;
            operation_274_2753 <= 32'd0;
            operation_274_2752 <= 32'd0;
            operation_274_2751 <= 32'd0;
            operation_274_2750 <= 32'd0;
            operation_274_2749 <= 32'd0;
            operation_274_2748 <= 32'd0;
            operation_274_2747 <= 32'd0;
            operation_274_2746 <= 32'd0;
            operation_274_2745 <= 32'd0;
            operation_274_2744 <= 32'd0;
            operation_274_2743 <= 32'd0;
            operation_274_2778 <= 32'd0;
            operation_274_2777 <= 32'd0;
            operation_274_2776 <= 32'd0;
            operation_274_2775 <= 32'd0;
            operation_274_2774 <= 32'd0;
            operation_274_2773 <= 32'd0;
            operation_274_2772 <= 32'd0;
            operation_274_2771 <= 32'd0;
            operation_274_2770 <= 32'd0;
            operation_274_2769 <= 32'd0;
            operation_274_2768 <= 32'd0;
            operation_274_2767 <= 32'd0;
            operation_274_2766 <= 32'd0;
            operation_274_2765 <= 32'd0;
            operation_274_2764 <= 32'd0;
            operation_274_2763 <= 32'd0;
            operation_274_2802 <= 32'd0;
            operation_274_2801 <= 32'd0;
            operation_274_2800 <= 32'd0;
            operation_274_2799 <= 32'd0;
            operation_274_2798 <= 32'd0;
            operation_274_2797 <= 32'd0;
            operation_274_2796 <= 32'd0;
            operation_274_2795 <= 32'd0;
            operation_274_2794 <= 32'd0;
            operation_274_2793 <= 32'd0;
            operation_274_2792 <= 32'd0;
            operation_274_2791 <= 32'd0;
            operation_274_2790 <= 32'd0;
            operation_274_2789 <= 32'd0;
            operation_274_2788 <= 32'd0;
            operation_274_2787 <= 32'd0;
            operation_274_3273 <= 32'd0;
            operation_274_3272 <= 32'd0;
            operation_274_3234 <= 32'd0;
            operation_274_3171 <= 32'd0;
            operation_274_2840 <= 32'd0;
            operation_274_2839 <= 32'd0;
            operation_274_2838 <= 32'd0;
            operation_274_2837 <= 32'd0;
            operation_274_2836 <= 32'd0;
            operation_274_2835 <= 32'd0;
            operation_274_2834 <= 32'd0;
            operation_274_2833 <= 32'd0;
            operation_274_2832 <= 32'd0;
            operation_274_2831 <= 32'd0;
            operation_274_2830 <= 32'd0;
            operation_274_2829 <= 32'd0;
            operation_274_2828 <= 32'd0;
            operation_274_2827 <= 32'd0;
            operation_274_2826 <= 32'd0;
            operation_274_2825 <= 32'd0;
            operation_274_2824 <= 32'd0;
            operation_274_2823 <= 32'd0;
            operation_274_2822 <= 32'd0;
            operation_274_2821 <= 32'd0;
            operation_274_2820 <= 32'd0;
            operation_274_2819 <= 32'd0;
            operation_274_2818 <= 32'd0;
            operation_274_2817 <= 32'd0;
            operation_274_2816 <= 32'd0;
            operation_274_2815 <= 32'd0;
            operation_274_2814 <= 32'd0;
            operation_274_2813 <= 32'd0;
            operation_274_2812 <= 32'd0;
            operation_274_2811 <= 32'd0;
            operation_274_2810 <= 32'd0;
            operation_274_2809 <= 32'd0;
            operation_274_2866 <= 32'd0;
            operation_274_2865 <= 32'd0;
            operation_274_2848 <= 32'd0;
            operation_274_2847 <= 32'd0;
            operation_274_2890 <= 32'd0;
            operation_274_2889 <= 32'd0;
            operation_274_2872 <= 32'd0;
            operation_274_2871 <= 32'd0;
            operation_274_3343 <= 32'd0;
            operation_274_3342 <= 32'd0;
            operation_274_3324 <= 32'd0;
            operation_274_3235 <= 32'd0;
            operation_274_2911 <= 32'd0;
            operation_274_2910 <= 32'd0;
            operation_274_2909 <= 32'd0;
            operation_274_2908 <= 32'd0;
            operation_274_2907 <= 32'd0;
            operation_274_2906 <= 32'd0;
            operation_274_2905 <= 32'd0;
            operation_274_2904 <= 32'd0;
            operation_274_2903 <= 32'd0;
            operation_274_2902 <= 32'd0;
            operation_274_2901 <= 32'd0;
            operation_274_2900 <= 32'd0;
            operation_274_2899 <= 32'd0;
            operation_274_2898 <= 32'd0;
            operation_274_2897 <= 32'd0;
            operation_274_2896 <= 32'd0;
            operation_274_3393_latch <= 8'd0;
            operation_274_3375_latch <= 8'd0;
            operation_274_3374_latch <= 8'd0;
            operation_274_2962_latch <= 8'd0;
            operation_274_2961_latch <= 8'd0;
            operation_274_2960_latch <= 8'd0;
            operation_274_2959_latch <= 8'd0;
            operation_274_2958_latch <= 8'd0;
            operation_274_2957_latch <= 8'd0;
            operation_274_2956_latch <= 8'd0;
            operation_274_2955_latch <= 8'd0;
            operation_274_2954_latch <= 8'd0;
            operation_274_2953_latch <= 8'd0;
            operation_274_2952_latch <= 8'd0;
            operation_274_2951_latch <= 8'd0;
            operation_274_2950_latch <= 8'd0;
            operation_274_2949_latch <= 8'd0;
            operation_274_2948_latch <= 8'd0;
            operation_274_2947_latch <= 8'd0;
            operation_274_3341 <= 32'd0;
            operation_274_2700 <= 32'd0;
            operation_274_2681 <= 32'd0;
            operation_274_2624 <= 32'd0;
            operation_274_2159 <= 32'd0;
            operation_274_2158 <= 32'd0;
            operation_274_2157 <= 32'd0;
            operation_274_2156 <= 32'd0;
            operation_274_2155 <= 32'd0;
            operation_274_2154 <= 32'd0;
            operation_274_2153 <= 32'd0;
            operation_274_2152 <= 32'd0;
            operation_274_2151 <= 32'd0;
            operation_274_2150 <= 32'd0;
            operation_274_2149 <= 32'd0;
            operation_274_2148 <= 32'd0;
            operation_274_2147 <= 32'd0;
            operation_274_2146 <= 32'd0;
            operation_274_2145 <= 32'd0;
            operation_274_2144 <= 32'd0;
            operation_274_3392_latch <= 8'd0;
            operation_274_2760 <= 32'd0;
            operation_274_2741 <= 32'd0;
            operation_274_2699 <= 32'd0;
            operation_274_2682 <= 32'd0;
            operation_274_2211 <= 32'd0;
            operation_274_2210 <= 32'd0;
            operation_274_2209 <= 32'd0;
            operation_274_2208 <= 32'd0;
            operation_274_2207 <= 32'd0;
            operation_274_2206 <= 32'd0;
            operation_274_2205 <= 32'd0;
            operation_274_2204 <= 32'd0;
            operation_274_2203 <= 32'd0;
            operation_274_2202 <= 32'd0;
            operation_274_2201 <= 32'd0;
            operation_274_2200 <= 32'd0;
            operation_274_2199 <= 32'd0;
            operation_274_2198 <= 32'd0;
            operation_274_2197 <= 32'd0;
            operation_274_2196 <= 32'd0;
            operation_274_2844 <= 32'd0;
            operation_274_2805 <= 32'd0;
            operation_274_2759 <= 32'd0;
            operation_274_2742 <= 32'd0;
            operation_274_2269 <= 32'd0;
            operation_274_2268 <= 32'd0;
            operation_274_2267 <= 32'd0;
            operation_274_2266 <= 32'd0;
            operation_274_2265 <= 32'd0;
            operation_274_2264 <= 32'd0;
            operation_274_2263 <= 32'd0;
            operation_274_2262 <= 32'd0;
            operation_274_2261 <= 32'd0;
            operation_274_2260 <= 32'd0;
            operation_274_2259 <= 32'd0;
            operation_274_2258 <= 32'd0;
            operation_274_2257 <= 32'd0;
            operation_274_2256 <= 32'd0;
            operation_274_2255 <= 32'd0;
            operation_274_2254 <= 32'd0;
            operation_274_2914 <= 32'd0;
            operation_274_2895 <= 32'd0;
            operation_274_2843 <= 32'd0;
            operation_274_2806 <= 32'd0;
            operation_274_2329 <= 32'd0;
            operation_274_2328 <= 32'd0;
            operation_274_2327 <= 32'd0;
            operation_274_2326 <= 32'd0;
            operation_274_2325 <= 32'd0;
            operation_274_2324 <= 32'd0;
            operation_274_2323 <= 32'd0;
            operation_274_2322 <= 32'd0;
            operation_274_2321 <= 32'd0;
            operation_274_2320 <= 32'd0;
            operation_274_2319 <= 32'd0;
            operation_274_2318 <= 32'd0;
            operation_274_2317 <= 32'd0;
            operation_274_2316 <= 32'd0;
            operation_274_2315 <= 32'd0;
            operation_274_2314 <= 32'd0;
            operation_274_2349 <= 32'd0;
            operation_274_2348 <= 32'd0;
            operation_274_2347 <= 32'd0;
            operation_274_2346 <= 32'd0;
            operation_274_2345 <= 32'd0;
            operation_274_2344 <= 32'd0;
            operation_274_2343 <= 32'd0;
            operation_274_2342 <= 32'd0;
            operation_274_2341 <= 32'd0;
            operation_274_2340 <= 32'd0;
            operation_274_2339 <= 32'd0;
            operation_274_2338 <= 32'd0;
            operation_274_2337 <= 32'd0;
            operation_274_2336 <= 32'd0;
            operation_274_2335 <= 32'd0;
            operation_274_2334 <= 32'd0;
            operation_274_2964_latch <= 8'd0;
            operation_274_2945_latch <= 8'd0;
            operation_274_2373 <= 32'd0;
            operation_274_2372 <= 32'd0;
            operation_274_2371 <= 32'd0;
            operation_274_2370 <= 32'd0;
            operation_274_2369 <= 32'd0;
            operation_274_2368 <= 32'd0;
            operation_274_2367 <= 32'd0;
            operation_274_2366 <= 32'd0;
            operation_274_2365 <= 32'd0;
            operation_274_2364 <= 32'd0;
            operation_274_2363 <= 32'd0;
            operation_274_2362 <= 32'd0;
            operation_274_2361 <= 32'd0;
            operation_274_2360 <= 32'd0;
            operation_274_2359 <= 32'd0;
            operation_274_2358 <= 32'd0;
            operation_274_2913 <= 32'd0;
            operation_274_2912 <= 32'd0;
            operation_274_2411 <= 32'd0;
            operation_274_2410 <= 32'd0;
            operation_274_2409 <= 32'd0;
            operation_274_2408 <= 32'd0;
            operation_274_2407 <= 32'd0;
            operation_274_2406 <= 32'd0;
            operation_274_2405 <= 32'd0;
            operation_274_2404 <= 32'd0;
            operation_274_2403 <= 32'd0;
            operation_274_2402 <= 32'd0;
            operation_274_2401 <= 32'd0;
            operation_274_2400 <= 32'd0;
            operation_274_2399 <= 32'd0;
            operation_274_2398 <= 32'd0;
            operation_274_2397 <= 32'd0;
            operation_274_2396 <= 32'd0;
            operation_274_2395 <= 32'd0;
            operation_274_2394 <= 32'd0;
            operation_274_2393 <= 32'd0;
            operation_274_2392 <= 32'd0;
            operation_274_2391 <= 32'd0;
            operation_274_2390 <= 32'd0;
            operation_274_2389 <= 32'd0;
            operation_274_2388 <= 32'd0;
            operation_274_2387 <= 32'd0;
            operation_274_2386 <= 32'd0;
            operation_274_2385 <= 32'd0;
            operation_274_2384 <= 32'd0;
            operation_274_2383 <= 32'd0;
            operation_274_2382 <= 32'd0;
            operation_274_2381 <= 32'd0;
            operation_274_2380 <= 32'd0;
            operation_274_2271 <= 32'd0;
            operation_274_2195 <= 32'd0;
            operation_274_2437 <= 32'd0;
            operation_274_2436 <= 32'd0;
            operation_274_2419 <= 32'd0;
            operation_274_2418 <= 32'd0;
            operation_274_2963_latch <= 8'd0;
            operation_274_2946_latch <= 8'd0;
            operation_274_2461 <= 32'd0;
            operation_274_2460 <= 32'd0;
            operation_274_2443 <= 32'd0;
            operation_274_2442 <= 32'd0;
            operation_274_2482 <= 32'd0;
            operation_274_2481 <= 32'd0;
            operation_274_2480 <= 32'd0;
            operation_274_2479 <= 32'd0;
            operation_274_2478 <= 32'd0;
            operation_274_2477 <= 32'd0;
            operation_274_2476 <= 32'd0;
            operation_274_2475 <= 32'd0;
            operation_274_2474 <= 32'd0;
            operation_274_2473 <= 32'd0;
            operation_274_2472 <= 32'd0;
            operation_274_2471 <= 32'd0;
            operation_274_2470 <= 32'd0;
            operation_274_2469 <= 32'd0;
            operation_274_2468 <= 32'd0;
            operation_274_2467 <= 32'd0;
            operation_274_2331 <= 32'd0;
            operation_274_2270 <= 32'd0;
            operation_274_2253 <= 32'd0;
            operation_274_2252 <= 32'd0;
            operation_274_2533_latch <= 8'd0;
            operation_274_2532_latch <= 8'd0;
            operation_274_2531_latch <= 8'd0;
            operation_274_2530_latch <= 8'd0;
            operation_274_2529_latch <= 8'd0;
            operation_274_2528_latch <= 8'd0;
            operation_274_2527_latch <= 8'd0;
            operation_274_2526_latch <= 8'd0;
            operation_274_2525_latch <= 8'd0;
            operation_274_2524_latch <= 8'd0;
            operation_274_2523_latch <= 8'd0;
            operation_274_2522_latch <= 8'd0;
            operation_274_2521_latch <= 8'd0;
            operation_274_2520_latch <= 8'd0;
            operation_274_2519_latch <= 8'd0;
            operation_274_2518_latch <= 8'd0;
            operation_274_2415 <= 32'd0;
            operation_274_2330 <= 32'd0;
            operation_274_2313 <= 32'd0;
            operation_274_2312 <= 32'd0;
            operation_274_1730 <= 32'd0;
            operation_274_1729 <= 32'd0;
            operation_274_1728 <= 32'd0;
            operation_274_1727 <= 32'd0;
            operation_274_1726 <= 32'd0;
            operation_274_1725 <= 32'd0;
            operation_274_1724 <= 32'd0;
            operation_274_1723 <= 32'd0;
            operation_274_1722 <= 32'd0;
            operation_274_1721 <= 32'd0;
            operation_274_1720 <= 32'd0;
            operation_274_1719 <= 32'd0;
            operation_274_1718 <= 32'd0;
            operation_274_1717 <= 32'd0;
            operation_274_1716 <= 32'd0;
            operation_274_1715 <= 32'd0;
            operation_274_2485 <= 32'd0;
            operation_274_2414 <= 32'd0;
            operation_274_2377 <= 32'd0;
            operation_274_2376 <= 32'd0;
            operation_274_1782 <= 32'd0;
            operation_274_1781 <= 32'd0;
            operation_274_1780 <= 32'd0;
            operation_274_1779 <= 32'd0;
            operation_274_1778 <= 32'd0;
            operation_274_1777 <= 32'd0;
            operation_274_1776 <= 32'd0;
            operation_274_1775 <= 32'd0;
            operation_274_1774 <= 32'd0;
            operation_274_1773 <= 32'd0;
            operation_274_1772 <= 32'd0;
            operation_274_1771 <= 32'd0;
            operation_274_1770 <= 32'd0;
            operation_274_1769 <= 32'd0;
            operation_274_1768 <= 32'd0;
            operation_274_1767 <= 32'd0;
            operation_274_2516_latch <= 8'd0;
            operation_274_2484 <= 32'd0;
            operation_274_2483 <= 32'd0;
            operation_274_2466 <= 32'd0;
            operation_274_1840 <= 32'd0;
            operation_274_1839 <= 32'd0;
            operation_274_1838 <= 32'd0;
            operation_274_1837 <= 32'd0;
            operation_274_1836 <= 32'd0;
            operation_274_1835 <= 32'd0;
            operation_274_1834 <= 32'd0;
            operation_274_1833 <= 32'd0;
            operation_274_1832 <= 32'd0;
            operation_274_1831 <= 32'd0;
            operation_274_1830 <= 32'd0;
            operation_274_1829 <= 32'd0;
            operation_274_1828 <= 32'd0;
            operation_274_1827 <= 32'd0;
            operation_274_1826 <= 32'd0;
            operation_274_1825 <= 32'd0;
            operation_274_1766 <= 32'd0;
            operation_274_2535_latch <= 8'd0;
            operation_274_2534_latch <= 8'd0;
            operation_274_2517_latch <= 8'd0;
            operation_274_1900 <= 32'd0;
            operation_274_1899 <= 32'd0;
            operation_274_1898 <= 32'd0;
            operation_274_1897 <= 32'd0;
            operation_274_1896 <= 32'd0;
            operation_274_1895 <= 32'd0;
            operation_274_1894 <= 32'd0;
            operation_274_1893 <= 32'd0;
            operation_274_1892 <= 32'd0;
            operation_274_1891 <= 32'd0;
            operation_274_1890 <= 32'd0;
            operation_274_1889 <= 32'd0;
            operation_274_1888 <= 32'd0;
            operation_274_1887 <= 32'd0;
            operation_274_1886 <= 32'd0;
            operation_274_1885 <= 32'd0;
            operation_274_1842 <= 32'd0;
            operation_274_1841 <= 32'd0;
            operation_274_1824 <= 32'd0;
            operation_274_1823 <= 32'd0;
            operation_274_1920 <= 32'd0;
            operation_274_1919 <= 32'd0;
            operation_274_1918 <= 32'd0;
            operation_274_1917 <= 32'd0;
            operation_274_1916 <= 32'd0;
            operation_274_1915 <= 32'd0;
            operation_274_1914 <= 32'd0;
            operation_274_1913 <= 32'd0;
            operation_274_1912 <= 32'd0;
            operation_274_1911 <= 32'd0;
            operation_274_1910 <= 32'd0;
            operation_274_1909 <= 32'd0;
            operation_274_1908 <= 32'd0;
            operation_274_1907 <= 32'd0;
            operation_274_1906 <= 32'd0;
            operation_274_1905 <= 32'd0;
            operation_274_1944 <= 32'd0;
            operation_274_1943 <= 32'd0;
            operation_274_1942 <= 32'd0;
            operation_274_1941 <= 32'd0;
            operation_274_1940 <= 32'd0;
            operation_274_1939 <= 32'd0;
            operation_274_1938 <= 32'd0;
            operation_274_1937 <= 32'd0;
            operation_274_1936 <= 32'd0;
            operation_274_1935 <= 32'd0;
            operation_274_1934 <= 32'd0;
            operation_274_1933 <= 32'd0;
            operation_274_1932 <= 32'd0;
            operation_274_1931 <= 32'd0;
            operation_274_1930 <= 32'd0;
            operation_274_1929 <= 32'd0;
            operation_274_1982 <= 32'd0;
            operation_274_1981 <= 32'd0;
            operation_274_1980 <= 32'd0;
            operation_274_1979 <= 32'd0;
            operation_274_1978 <= 32'd0;
            operation_274_1977 <= 32'd0;
            operation_274_1976 <= 32'd0;
            operation_274_1975 <= 32'd0;
            operation_274_1974 <= 32'd0;
            operation_274_1973 <= 32'd0;
            operation_274_1972 <= 32'd0;
            operation_274_1971 <= 32'd0;
            operation_274_1970 <= 32'd0;
            operation_274_1969 <= 32'd0;
            operation_274_1968 <= 32'd0;
            operation_274_1967 <= 32'd0;
            operation_274_1966 <= 32'd0;
            operation_274_1965 <= 32'd0;
            operation_274_1964 <= 32'd0;
            operation_274_1963 <= 32'd0;
            operation_274_1962 <= 32'd0;
            operation_274_1961 <= 32'd0;
            operation_274_1960 <= 32'd0;
            operation_274_1959 <= 32'd0;
            operation_274_1958 <= 32'd0;
            operation_274_1957 <= 32'd0;
            operation_274_1956 <= 32'd0;
            operation_274_1955 <= 32'd0;
            operation_274_1954 <= 32'd0;
            operation_274_1953 <= 32'd0;
            operation_274_1952 <= 32'd0;
            operation_274_1951 <= 32'd0;
            operation_274_1902 <= 32'd0;
            operation_274_1901 <= 32'd0;
            operation_274_1884 <= 32'd0;
            operation_274_1883 <= 32'd0;
            operation_274_2008 <= 32'd0;
            operation_274_2007 <= 32'd0;
            operation_274_1990 <= 32'd0;
            operation_274_1989 <= 32'd0;
            operation_274_2032 <= 32'd0;
            operation_274_2031 <= 32'd0;
            operation_274_2014 <= 32'd0;
            operation_274_2013 <= 32'd0;
            operation_274_2053 <= 32'd0;
            operation_274_2052 <= 32'd0;
            operation_274_2051 <= 32'd0;
            operation_274_2050 <= 32'd0;
            operation_274_2049 <= 32'd0;
            operation_274_2048 <= 32'd0;
            operation_274_2047 <= 32'd0;
            operation_274_2046 <= 32'd0;
            operation_274_2045 <= 32'd0;
            operation_274_2044 <= 32'd0;
            operation_274_2043 <= 32'd0;
            operation_274_2042 <= 32'd0;
            operation_274_2041 <= 32'd0;
            operation_274_2040 <= 32'd0;
            operation_274_2039 <= 32'd0;
            operation_274_2038 <= 32'd0;
            operation_274_1986 <= 32'd0;
            operation_274_1985 <= 32'd0;
            operation_274_1948 <= 32'd0;
            operation_274_1947 <= 32'd0;
            operation_274_2104_latch <= 8'd0;
            operation_274_2103_latch <= 8'd0;
            operation_274_2102_latch <= 8'd0;
            operation_274_2101_latch <= 8'd0;
            operation_274_2100_latch <= 8'd0;
            operation_274_2099_latch <= 8'd0;
            operation_274_2098_latch <= 8'd0;
            operation_274_2097_latch <= 8'd0;
            operation_274_2096_latch <= 8'd0;
            operation_274_2095_latch <= 8'd0;
            operation_274_2094_latch <= 8'd0;
            operation_274_2093_latch <= 8'd0;
            operation_274_2092_latch <= 8'd0;
            operation_274_2091_latch <= 8'd0;
            operation_274_2090_latch <= 8'd0;
            operation_274_2089_latch <= 8'd0;
            operation_274_2056 <= 32'd0;
            operation_274_2055 <= 32'd0;
            operation_274_2054 <= 32'd0;
            operation_274_2037 <= 32'd0;
            operation_274_118 <= 32'd0;
            operation_274_102 <= 32'd0;
            operation_274_86 <= 32'd0;
            operation_274_70 <= 32'd0;
            operation_274_54 <= 32'd0;
            operation_274_38 <= 32'd0;
            operation_274_22 <= 32'd0;
            operation_274_6 <= 32'd0;
            operation_274_14 <= 32'd0;
            operation_274_30 <= 32'd0;
            operation_274_46 <= 32'd0;
            operation_274_62 <= 32'd0;
            operation_274_78 <= 32'd0;
            operation_274_94 <= 32'd0;
            operation_274_110 <= 32'd0;
            operation_274_126 <= 32'd0;
            operation_274_2106_latch <= 8'd0;
            operation_274_2105_latch <= 8'd0;
            operation_274_2088_latch <= 8'd0;
            operation_274_2087_latch <= 8'd0;
            control_274_follow <= 1'd0;
            control_274_start <= 1'd0;
            control_274_84 <= 1'd0;
            control_274_83 <= 1'd0;
            control_274_82 <= 1'd0;
            control_274_81 <= 1'd0;
            control_274_80 <= 1'd0;
            control_274_79 <= 1'd0;
            control_274_78 <= 1'd0;
            control_274_77 <= 1'd0;
            control_274_76 <= 1'd0;
            control_274_75 <= 1'd0;
            control_274_74 <= 1'd0;
            control_274_73 <= 1'd0;
            control_274_72 <= 1'd0;
            control_274_71 <= 1'd0;
            control_274_70 <= 1'd0;
            control_274_69 <= 1'd0;
            control_274_68 <= 1'd0;
            control_274_67 <= 1'd0;
            control_274_66 <= 1'd0;
            control_274_65 <= 1'd0;
            control_274_64 <= 1'd0;
            control_274_63 <= 1'd0;
            control_274_62 <= 1'd0;
            control_274_61 <= 1'd0;
            control_274_60 <= 1'd0;
            control_274_59 <= 1'd0;
            control_274_58 <= 1'd0;
            control_274_57 <= 1'd0;
            control_274_56 <= 1'd0;
            control_274_55 <= 1'd0;
            control_274_54 <= 1'd0;
            control_274_53 <= 1'd0;
            control_274_52 <= 1'd0;
            control_274_51 <= 1'd0;
            control_274_50 <= 1'd0;
            control_274_49 <= 1'd0;
            control_274_48 <= 1'd0;
            control_274_47 <= 1'd0;
            control_274_46 <= 1'd0;
            control_274_45 <= 1'd0;
            control_274_44 <= 1'd0;
            control_274_43 <= 1'd0;
            control_274_42 <= 1'd0;
            control_274_41 <= 1'd0;
            control_274_40 <= 1'd0;
            control_274_39 <= 1'd0;
            control_274_38 <= 1'd0;
            control_274_37 <= 1'd0;
            control_274_36 <= 1'd0;
            control_274_35 <= 1'd0;
            control_274_34 <= 1'd0;
            control_274_33 <= 1'd0;
            control_274_32 <= 1'd0;
            control_274_31 <= 1'd0;
            control_274_30 <= 1'd0;
            control_274_29 <= 1'd0;
            control_274_28 <= 1'd0;
            control_274_27 <= 1'd0;
            control_274_26 <= 1'd0;
            control_274_25 <= 1'd0;
            control_274_24 <= 1'd0;
            control_274_23 <= 1'd0;
            control_274_22 <= 1'd0;
            control_274_21 <= 1'd0;
            control_274_20 <= 1'd0;
            control_274_19 <= 1'd0;
            control_274_18 <= 1'd0;
            control_274_17 <= 1'd0;
            control_274_16 <= 1'd0;
            control_274_15 <= 1'd0;
            control_274_14 <= 1'd0;
            control_274_13 <= 1'd0;
            control_274_12 <= 1'd0;
            control_274_11 <= 1'd0;
            control_274_10 <= 1'd0;
            control_274_9 <= 1'd0;
            control_274_8 <= 1'd0;
            control_274_7 <= 1'd0;
            control_274_6 <= 1'd0;
            control_274_5 <= 1'd0;
            control_274_4 <= 1'd0;
            control_274_3 <= 1'd0;
            control_274_2 <= 1'd0;
            control_274_1 <= 1'd0;
            input_key_274_follow <= 128'd0;
            input_in_274_follow <= 128'd0;
            lookup_sbox_0_output <= 8'd0;
            lookup_sbox_1_output <= 8'd0;
            lookup_sbox_2_output <= 8'd0;
            lookup_sbox_3_output <= 8'd0;
            lookup_sbox_4_output <= 8'd0;
            lookup_sbox_5_output <= 8'd0;
            lookup_sbox_6_output <= 8'd0;
            lookup_sbox_7_output <= 8'd0;
            lookup_sbox_8_output <= 8'd0;
            lookup_sbox_9_output <= 8'd0;
            lookup_sbox_10_output <= 8'd0;
            lookup_sbox_11_output <= 8'd0;
            lookup_sbox_12_output <= 8'd0;
            lookup_sbox_13_output <= 8'd0;
            lookup_sbox_14_output <= 8'd0;
            lookup_sbox_15_output <= 8'd0;
            startfollow <= 1'd0;
        end
    else
        begin
            AES128_encrypt <= ((control_274_follow)?(return_274):(AES128_encrypt));
            finish <= (((finish)&&(!((start)&&(!(startfollow)))))||(control_274_end));
            control_274_start <= ((start)&&(!(startfollow)));
            operation_274_1664 <= ((operation_274_1661)^(operation_274_1663));
            operation_274_1688 <= ((operation_274_1685)^(operation_274_1687));
            operation_274_1672 <= ((operation_274_1669)^(operation_274_1671));
            operation_274_1632 <= ((operation_274_1629)^(operation_274_1535));
            operation_274_1680 <= ((operation_274_1677)^(operation_274_1679));
            operation_274_1656 <= ((operation_274_1653)^(operation_274_1655));
            operation_274_1640 <= ((operation_274_1637)^(operation_274_1639));
            operation_274_1600 <= ((operation_274_1597)^(operation_274_1503));
            operation_274_1648 <= ((operation_274_1645)^(operation_274_1551));
            operation_274_1624 <= ((operation_274_1621)^(operation_274_1623));
            operation_274_1608 <= ((operation_274_1605)^(operation_274_1607));
            operation_274_1568 <= ((operation_274_1565)^(operation_274_1471));
            operation_274_1616 <= ((operation_274_1613)^(operation_274_1519));
            operation_274_1592 <= ((operation_274_1589)^(operation_274_1591));
            operation_274_1576 <= ((operation_274_1573)^(operation_274_1575));
            operation_274_1584 <= ((operation_274_1581)^(operation_274_1487));
            operation_274_1338_latch <= (operation_274_1338);
            operation_274_1328_latch <= (operation_274_1328);
            operation_274_1318_latch <= (operation_274_1318);
            operation_274_1308_latch <= (operation_274_1308);
            operation_274_1298_latch <= (operation_274_1298);
            operation_274_1288_latch <= (operation_274_1288);
            operation_274_1278_latch <= (operation_274_1278);
            operation_274_1268_latch <= (operation_274_1268);
            operation_274_1273_latch <= (operation_274_1273);
            operation_274_1283_latch <= (operation_274_1283);
            operation_274_1293_latch <= (operation_274_1293);
            operation_274_1303_latch <= (operation_274_1303);
            operation_274_1313_latch <= (operation_274_1313);
            operation_274_1323_latch <= (operation_274_1323);
            operation_274_1333_latch <= (operation_274_1333);
            operation_274_1343_latch <= (operation_274_1343);
            operation_274_5162 <= ((operation_274_5180)^(operation_274_5234));
            operation_274_5161 <= ((operation_274_5179)^(operation_274_5233));
            operation_274_5160 <= ((operation_274_5178)^(operation_274_5294));
            operation_274_5159 <= ((operation_274_5177)^(operation_274_5293));
            operation_274_5158 <= ((operation_274_5176)^(operation_274_5354));
            operation_274_5157 <= ((operation_274_5175)^(operation_274_5353));
            operation_274_5156 <= ((operation_274_5174)^(operation_274_5442));
            operation_274_5155 <= ((operation_274_5173)^(operation_274_5441));
            operation_274_5154 <= ((operation_274_5171)^(operation_274_5336));
            operation_274_5153 <= ((operation_274_5170)^(operation_274_5419));
            operation_274_5152 <= ((operation_274_5169)^(operation_274_5276));
            operation_274_5151 <= ((operation_274_5168)^(operation_274_5335));
            operation_274_5150 <= ((operation_274_5167)^(operation_274_5216));
            operation_274_5149 <= ((operation_274_5166)^(operation_274_5275));
            operation_274_5148 <= ((operation_274_5165)^(operation_274_5164));
            operation_274_5147 <= ((operation_274_5163)^(operation_274_5215));
            operation_274_5214 <= ((operation_274_5501)^(operation_274_5232));
            operation_274_5213 <= ((operation_274_5500)^(operation_274_5231));
            operation_274_5212 <= ((operation_274_5505)^(operation_274_5230));
            operation_274_5211 <= ((operation_274_5504)^(operation_274_5229));
            operation_274_5210 <= ((operation_274_5503)^(operation_274_5228));
            operation_274_5209 <= ((operation_274_5502)^(operation_274_5227));
            operation_274_5208 <= ((operation_274_5507)^(operation_274_5226));
            operation_274_5207 <= ((operation_274_5506)^(operation_274_5225));
            operation_274_5206 <= ((operation_274_5499)^(operation_274_5224));
            operation_274_5205 <= ((operation_274_5498)^(operation_274_5223));
            operation_274_5204 <= ((operation_274_5497)^(operation_274_5222));
            operation_274_5203 <= ((operation_274_5496)^(operation_274_5221));
            operation_274_5202 <= ((operation_274_5495)^(operation_274_5220));
            operation_274_5201 <= ((operation_274_5494)^(operation_274_5219));
            operation_274_5200 <= ((operation_274_5493)^(operation_274_5218));
            operation_274_5199 <= ((operation_274_5492)^(operation_274_5217));
            operation_274_5272 <= ((operation_274_5292)^(operation_274_5357));
            operation_274_5271 <= ((operation_274_5291)^(operation_274_5357));
            operation_274_5270 <= ((operation_274_5290)^(operation_274_5358));
            operation_274_5269 <= ((operation_274_5289)^(operation_274_5358));
            operation_274_5268 <= ((operation_274_5288)^(operation_274_5359));
            operation_274_5267 <= ((operation_274_5287)^(operation_274_5359));
            operation_274_5266 <= ((operation_274_5286)^(operation_274_5360));
            operation_274_5265 <= ((operation_274_5285)^(operation_274_5360));
            operation_274_5264 <= ((operation_274_5284)^(operation_274_5360));
            operation_274_5263 <= ((operation_274_5283)^(operation_274_5360));
            operation_274_5262 <= ((operation_274_5282)^(operation_274_5359));
            operation_274_5261 <= ((operation_274_5281)^(operation_274_5359));
            operation_274_5260 <= ((operation_274_5280)^(operation_274_5358));
            operation_274_5259 <= ((operation_274_5279)^(operation_274_5358));
            operation_274_5258 <= ((operation_274_5278)^(operation_274_5357));
            operation_274_5257 <= ((operation_274_5277)^(operation_274_5357));
            operation_274_5332 <= ((operation_274_5413)^(operation_274_5352));
            operation_274_5331 <= ((operation_274_5411)^(operation_274_5351));
            operation_274_5330 <= ((operation_274_5409)^(operation_274_5350));
            operation_274_5329 <= ((operation_274_5407)^(operation_274_5349));
            operation_274_5328 <= ((operation_274_5405)^(operation_274_5348));
            operation_274_5327 <= ((operation_274_5403)^(operation_274_5347));
            operation_274_5326 <= ((operation_274_5401)^(operation_274_5346));
            operation_274_5325 <= ((operation_274_5399)^(operation_274_5345));
            operation_274_5324 <= ((operation_274_5398)^(operation_274_5344));
            operation_274_5323 <= ((operation_274_5396)^(operation_274_5343));
            operation_274_5322 <= ((operation_274_5394)^(operation_274_5342));
            operation_274_5321 <= ((operation_274_5392)^(operation_274_5341));
            operation_274_5320 <= ((operation_274_5390)^(operation_274_5340));
            operation_274_5319 <= ((operation_274_5388)^(operation_274_5339));
            operation_274_5318 <= ((operation_274_5386)^(operation_274_5338));
            operation_274_5317 <= ((operation_274_5384)^(operation_274_5337));
            operation_274_5352 <= ((operation_274_5376)*(operation_274_5597));
            operation_274_5351 <= ((operation_274_5375)*(operation_274_5597));
            operation_274_5350 <= ((operation_274_5374)*(operation_274_5597));
            operation_274_5349 <= ((operation_274_5373)*(operation_274_5597));
            operation_274_5348 <= ((operation_274_5372)*(operation_274_5597));
            operation_274_5347 <= ((operation_274_5371)*(operation_274_5597));
            operation_274_5346 <= ((operation_274_5370)*(operation_274_5597));
            operation_274_5345 <= ((operation_274_5369)*(operation_274_5597));
            operation_274_5344 <= ((operation_274_5368)*(operation_274_5597));
            operation_274_5343 <= ((operation_274_5367)*(operation_274_5597));
            operation_274_5342 <= ((operation_274_5366)*(operation_274_5597));
            operation_274_5341 <= ((operation_274_5365)*(operation_274_5597));
            operation_274_5340 <= ((operation_274_5364)*(operation_274_5597));
            operation_274_5339 <= ((operation_274_5363)*(operation_274_5597));
            operation_274_5338 <= ((operation_274_5362)*(operation_274_5597));
            operation_274_5337 <= ((operation_274_5361)*(operation_274_5597));
            operation_274_5376 <= ((operation_274_5414)&(operation_274_5557));
            operation_274_5375 <= ((operation_274_5412)&(operation_274_5557));
            operation_274_5374 <= ((operation_274_5410)&(operation_274_5557));
            operation_274_5373 <= ((operation_274_5408)&(operation_274_5557));
            operation_274_5372 <= ((operation_274_5406)&(operation_274_5557));
            operation_274_5371 <= ((operation_274_5404)&(operation_274_5557));
            operation_274_5370 <= ((operation_274_5402)&(operation_274_5557));
            operation_274_5369 <= ((operation_274_5400)&(operation_274_5557));
            operation_274_5368 <= ((operation_274_5397)&(operation_274_5557));
            operation_274_5367 <= ((operation_274_5395)&(operation_274_5557));
            operation_274_5366 <= ((operation_274_5393)&(operation_274_5557));
            operation_274_5365 <= ((operation_274_5391)&(operation_274_5557));
            operation_274_5364 <= ((operation_274_5389)&(operation_274_5557));
            operation_274_5363 <= ((operation_274_5387)&(operation_274_5557));
            operation_274_5362 <= ((operation_274_5385)&(operation_274_5557));
            operation_274_5361 <= ((operation_274_5383)&(operation_274_5557));
            operation_274_5414 <= ((operation_274_5438)>>(operation_274_2119));
            operation_274_5413 <= ((operation_274_5438)<<(operation_274_5557));
            operation_274_5412 <= ((operation_274_5437)>>(operation_274_2119));
            operation_274_5411 <= ((operation_274_5437)<<(operation_274_5557));
            operation_274_5410 <= ((operation_274_5436)>>(operation_274_2119));
            operation_274_5409 <= ((operation_274_5436)<<(operation_274_5557));
            operation_274_5408 <= ((operation_274_5435)>>(operation_274_2119));
            operation_274_5407 <= ((operation_274_5435)<<(operation_274_5557));
            operation_274_5406 <= ((operation_274_5434)>>(operation_274_2119));
            operation_274_5405 <= ((operation_274_5434)<<(operation_274_5557));
            operation_274_5404 <= ((operation_274_5433)>>(operation_274_2119));
            operation_274_5403 <= ((operation_274_5433)<<(operation_274_5557));
            operation_274_5402 <= ((operation_274_5432)>>(operation_274_2119));
            operation_274_5401 <= ((operation_274_5432)<<(operation_274_5557));
            operation_274_5400 <= ((operation_274_5431)>>(operation_274_2119));
            operation_274_5399 <= ((operation_274_5431)<<(operation_274_5557));
            operation_274_5398 <= ((operation_274_5430)<<(operation_274_5557));
            operation_274_5397 <= ((operation_274_5430)>>(operation_274_2119));
            operation_274_5396 <= ((operation_274_5429)<<(operation_274_5557));
            operation_274_5395 <= ((operation_274_5429)>>(operation_274_2119));
            operation_274_5394 <= ((operation_274_5428)<<(operation_274_5557));
            operation_274_5393 <= ((operation_274_5428)>>(operation_274_2119));
            operation_274_5392 <= ((operation_274_5427)<<(operation_274_5557));
            operation_274_5391 <= ((operation_274_5427)>>(operation_274_2119));
            operation_274_5390 <= ((operation_274_5426)<<(operation_274_5557));
            operation_274_5389 <= ((operation_274_5426)>>(operation_274_2119));
            operation_274_5388 <= ((operation_274_5425)<<(operation_274_5557));
            operation_274_5387 <= ((operation_274_5425)>>(operation_274_2119));
            operation_274_5386 <= ((operation_274_5424)<<(operation_274_5557));
            operation_274_5385 <= ((operation_274_5424)>>(operation_274_2119));
            operation_274_5384 <= ((operation_274_5423)<<(operation_274_5557));
            operation_274_5383 <= ((operation_274_5423)>>(operation_274_2119));
            operation_274_5440 <= ((operation_274_5464)^(operation_274_5494));
            operation_274_5439 <= ((operation_274_5463)^(operation_274_5498));
            operation_274_5422 <= ((operation_274_5446)^(operation_274_5496));
            operation_274_5421 <= ((operation_274_5445)^(operation_274_5492));
            operation_274_5464 <= ((operation_274_5483)^(operation_274_5505));
            operation_274_5463 <= ((operation_274_5480)^(operation_274_5507));
            operation_274_5446 <= ((operation_274_5471)^(operation_274_5503));
            operation_274_5445 <= ((operation_274_5470)^(operation_274_5501));
            operation_274_5485 <= ((operation_274_5501)^(operation_274_5492));
            operation_274_5484 <= ((operation_274_5505)^(operation_274_5494));
            operation_274_5483 <= ((operation_274_5504)^(operation_274_5495));
            operation_274_5482 <= ((operation_274_5503)^(operation_274_5496));
            operation_274_5481 <= ((operation_274_5507)^(operation_274_5498));
            operation_274_5480 <= ((operation_274_5506)^(operation_274_5499));
            operation_274_5479 <= ((operation_274_5499)^(operation_274_5507));
            operation_274_5478 <= ((operation_274_5498)^(operation_274_5506));
            operation_274_5477 <= ((operation_274_5497)^(operation_274_5503));
            operation_274_5476 <= ((operation_274_5496)^(operation_274_5502));
            operation_274_5475 <= ((operation_274_5495)^(operation_274_5505));
            operation_274_5474 <= ((operation_274_5494)^(operation_274_5504));
            operation_274_5473 <= ((operation_274_5493)^(operation_274_5501));
            operation_274_5472 <= ((operation_274_5492)^(operation_274_5500));
            operation_274_5471 <= ((operation_274_5502)^(operation_274_5497));
            operation_274_5470 <= ((operation_274_5500)^(operation_274_5493));
            operation_274_5536_latch <= (operation_274_5536);
            operation_274_5535_latch <= (operation_274_5535);
            operation_274_5534_latch <= (operation_274_5534);
            operation_274_5533_latch <= (operation_274_5533);
            operation_274_5532_latch <= (operation_274_5532);
            operation_274_5531_latch <= (operation_274_5531);
            operation_274_5530_latch <= (operation_274_5530);
            operation_274_5529_latch <= (operation_274_5529);
            operation_274_5528_latch <= (operation_274_5528);
            operation_274_5527_latch <= (operation_274_5527);
            operation_274_5526_latch <= (operation_274_5526);
            operation_274_5525_latch <= (operation_274_5525);
            operation_274_5524_latch <= (operation_274_5524);
            operation_274_5523_latch <= (operation_274_5523);
            operation_274_5522_latch <= (operation_274_5522);
            operation_274_5521_latch <= (operation_274_5521);
            operation_274_4733 <= ((operation_274_4751)^(operation_274_4805));
            operation_274_4732 <= ((operation_274_4750)^(operation_274_4804));
            operation_274_4731 <= ((operation_274_4749)^(operation_274_4865));
            operation_274_4730 <= ((operation_274_4748)^(operation_274_4864));
            operation_274_4729 <= ((operation_274_4747)^(operation_274_4925));
            operation_274_4728 <= ((operation_274_4746)^(operation_274_4924));
            operation_274_4727 <= ((operation_274_4745)^(operation_274_5013));
            operation_274_4726 <= ((operation_274_4744)^(operation_274_5012));
            operation_274_4725 <= ((operation_274_4742)^(operation_274_4907));
            operation_274_4724 <= ((operation_274_4741)^(operation_274_4990));
            operation_274_4723 <= ((operation_274_4740)^(operation_274_4847));
            operation_274_4722 <= ((operation_274_4739)^(operation_274_4906));
            operation_274_4721 <= ((operation_274_4738)^(operation_274_4787));
            operation_274_4720 <= ((operation_274_4737)^(operation_274_4846));
            operation_274_4719 <= ((operation_274_4736)^(operation_274_4735));
            operation_274_4718 <= ((operation_274_4734)^(operation_274_4786));
            operation_274_4785 <= ((operation_274_5072)^(operation_274_4803));
            operation_274_4784 <= ((operation_274_5071)^(operation_274_4802));
            operation_274_4783 <= ((operation_274_5076)^(operation_274_4801));
            operation_274_4782 <= ((operation_274_5075)^(operation_274_4800));
            operation_274_4781 <= ((operation_274_5074)^(operation_274_4799));
            operation_274_4780 <= ((operation_274_5073)^(operation_274_4798));
            operation_274_4779 <= ((operation_274_5078)^(operation_274_4797));
            operation_274_4778 <= ((operation_274_5077)^(operation_274_4796));
            operation_274_4777 <= ((operation_274_5070)^(operation_274_4795));
            operation_274_4776 <= ((operation_274_5069)^(operation_274_4794));
            operation_274_4775 <= ((operation_274_5068)^(operation_274_4793));
            operation_274_4774 <= ((operation_274_5067)^(operation_274_4792));
            operation_274_4773 <= ((operation_274_5066)^(operation_274_4791));
            operation_274_4772 <= ((operation_274_5065)^(operation_274_4790));
            operation_274_4771 <= ((operation_274_5064)^(operation_274_4789));
            operation_274_4770 <= ((operation_274_5063)^(operation_274_4788));
            operation_274_4843 <= ((operation_274_4863)^(operation_274_4928));
            operation_274_4842 <= ((operation_274_4862)^(operation_274_4928));
            operation_274_4841 <= ((operation_274_4861)^(operation_274_4929));
            operation_274_4840 <= ((operation_274_4860)^(operation_274_4929));
            operation_274_4839 <= ((operation_274_4859)^(operation_274_4930));
            operation_274_4838 <= ((operation_274_4858)^(operation_274_4930));
            operation_274_4837 <= ((operation_274_4857)^(operation_274_4931));
            operation_274_4836 <= ((operation_274_4856)^(operation_274_4931));
            operation_274_4835 <= ((operation_274_4855)^(operation_274_4931));
            operation_274_4834 <= ((operation_274_4854)^(operation_274_4931));
            operation_274_4833 <= ((operation_274_4853)^(operation_274_4930));
            operation_274_4832 <= ((operation_274_4852)^(operation_274_4930));
            operation_274_4831 <= ((operation_274_4851)^(operation_274_4929));
            operation_274_4830 <= ((operation_274_4850)^(operation_274_4929));
            operation_274_4829 <= ((operation_274_4849)^(operation_274_4928));
            operation_274_4828 <= ((operation_274_4848)^(operation_274_4928));
            operation_274_4903 <= ((operation_274_4984)^(operation_274_4923));
            operation_274_4902 <= ((operation_274_4982)^(operation_274_4922));
            operation_274_4901 <= ((operation_274_4980)^(operation_274_4921));
            operation_274_4900 <= ((operation_274_4978)^(operation_274_4920));
            operation_274_4899 <= ((operation_274_4976)^(operation_274_4919));
            operation_274_4898 <= ((operation_274_4974)^(operation_274_4918));
            operation_274_4897 <= ((operation_274_4972)^(operation_274_4917));
            operation_274_4896 <= ((operation_274_4970)^(operation_274_4916));
            operation_274_4895 <= ((operation_274_4969)^(operation_274_4915));
            operation_274_4894 <= ((operation_274_4967)^(operation_274_4914));
            operation_274_4893 <= ((operation_274_4965)^(operation_274_4913));
            operation_274_4892 <= ((operation_274_4963)^(operation_274_4912));
            operation_274_4891 <= ((operation_274_4961)^(operation_274_4911));
            operation_274_4890 <= ((operation_274_4959)^(operation_274_4910));
            operation_274_4889 <= ((operation_274_4957)^(operation_274_4909));
            operation_274_4888 <= ((operation_274_4955)^(operation_274_4908));
            operation_274_4923 <= ((operation_274_4947)*(operation_274_5597));
            operation_274_4922 <= ((operation_274_4946)*(operation_274_5597));
            operation_274_4921 <= ((operation_274_4945)*(operation_274_5597));
            operation_274_4920 <= ((operation_274_4944)*(operation_274_5597));
            operation_274_4919 <= ((operation_274_4943)*(operation_274_5597));
            operation_274_4918 <= ((operation_274_4942)*(operation_274_5597));
            operation_274_4917 <= ((operation_274_4941)*(operation_274_5597));
            operation_274_4916 <= ((operation_274_4940)*(operation_274_5597));
            operation_274_4915 <= ((operation_274_4939)*(operation_274_5597));
            operation_274_4914 <= ((operation_274_4938)*(operation_274_5597));
            operation_274_4913 <= ((operation_274_4937)*(operation_274_5597));
            operation_274_4912 <= ((operation_274_4936)*(operation_274_5597));
            operation_274_4911 <= ((operation_274_4935)*(operation_274_5597));
            operation_274_4910 <= ((operation_274_4934)*(operation_274_5597));
            operation_274_4909 <= ((operation_274_4933)*(operation_274_5597));
            operation_274_4908 <= ((operation_274_4932)*(operation_274_5597));
            operation_274_4947 <= ((operation_274_4985)&(operation_274_5557));
            operation_274_4946 <= ((operation_274_4983)&(operation_274_5557));
            operation_274_4945 <= ((operation_274_4981)&(operation_274_5557));
            operation_274_4944 <= ((operation_274_4979)&(operation_274_5557));
            operation_274_4943 <= ((operation_274_4977)&(operation_274_5557));
            operation_274_4942 <= ((operation_274_4975)&(operation_274_5557));
            operation_274_4941 <= ((operation_274_4973)&(operation_274_5557));
            operation_274_4940 <= ((operation_274_4971)&(operation_274_5557));
            operation_274_4939 <= ((operation_274_4968)&(operation_274_5557));
            operation_274_4938 <= ((operation_274_4966)&(operation_274_5557));
            operation_274_4937 <= ((operation_274_4964)&(operation_274_5557));
            operation_274_4936 <= ((operation_274_4962)&(operation_274_5557));
            operation_274_4935 <= ((operation_274_4960)&(operation_274_5557));
            operation_274_4934 <= ((operation_274_4958)&(operation_274_5557));
            operation_274_4933 <= ((operation_274_4956)&(operation_274_5557));
            operation_274_4932 <= ((operation_274_4954)&(operation_274_5557));
            operation_274_4985 <= ((operation_274_5009)>>(operation_274_2119));
            operation_274_4984 <= ((operation_274_5009)<<(operation_274_5557));
            operation_274_4983 <= ((operation_274_5008)>>(operation_274_2119));
            operation_274_4982 <= ((operation_274_5008)<<(operation_274_5557));
            operation_274_4981 <= ((operation_274_5007)>>(operation_274_2119));
            operation_274_4980 <= ((operation_274_5007)<<(operation_274_5557));
            operation_274_4979 <= ((operation_274_5006)>>(operation_274_2119));
            operation_274_4978 <= ((operation_274_5006)<<(operation_274_5557));
            operation_274_4977 <= ((operation_274_5005)>>(operation_274_2119));
            operation_274_4976 <= ((operation_274_5005)<<(operation_274_5557));
            operation_274_4975 <= ((operation_274_5004)>>(operation_274_2119));
            operation_274_4974 <= ((operation_274_5004)<<(operation_274_5557));
            operation_274_4973 <= ((operation_274_5003)>>(operation_274_2119));
            operation_274_4972 <= ((operation_274_5003)<<(operation_274_5557));
            operation_274_4971 <= ((operation_274_5002)>>(operation_274_2119));
            operation_274_4970 <= ((operation_274_5002)<<(operation_274_5557));
            operation_274_4969 <= ((operation_274_5001)<<(operation_274_5557));
            operation_274_4968 <= ((operation_274_5001)>>(operation_274_2119));
            operation_274_4967 <= ((operation_274_5000)<<(operation_274_5557));
            operation_274_4966 <= ((operation_274_5000)>>(operation_274_2119));
            operation_274_4965 <= ((operation_274_4999)<<(operation_274_5557));
            operation_274_4964 <= ((operation_274_4999)>>(operation_274_2119));
            operation_274_4963 <= ((operation_274_4998)<<(operation_274_5557));
            operation_274_4962 <= ((operation_274_4998)>>(operation_274_2119));
            operation_274_4961 <= ((operation_274_4997)<<(operation_274_5557));
            operation_274_4960 <= ((operation_274_4997)>>(operation_274_2119));
            operation_274_4959 <= ((operation_274_4996)<<(operation_274_5557));
            operation_274_4958 <= ((operation_274_4996)>>(operation_274_2119));
            operation_274_4957 <= ((operation_274_4995)<<(operation_274_5557));
            operation_274_4956 <= ((operation_274_4995)>>(operation_274_2119));
            operation_274_4955 <= ((operation_274_4994)<<(operation_274_5557));
            operation_274_4954 <= ((operation_274_4994)>>(operation_274_2119));
            operation_274_5011 <= ((operation_274_5035)^(operation_274_5065));
            operation_274_5010 <= ((operation_274_5034)^(operation_274_5069));
            operation_274_4993 <= ((operation_274_5017)^(operation_274_5067));
            operation_274_4992 <= ((operation_274_5016)^(operation_274_5063));
            operation_274_5035 <= ((operation_274_5054)^(operation_274_5076));
            operation_274_5034 <= ((operation_274_5051)^(operation_274_5078));
            operation_274_5017 <= ((operation_274_5042)^(operation_274_5074));
            operation_274_5016 <= ((operation_274_5041)^(operation_274_5072));
            operation_274_5056 <= ((operation_274_5072)^(operation_274_5063));
            operation_274_5055 <= ((operation_274_5076)^(operation_274_5065));
            operation_274_5054 <= ((operation_274_5075)^(operation_274_5066));
            operation_274_5053 <= ((operation_274_5074)^(operation_274_5067));
            operation_274_5052 <= ((operation_274_5078)^(operation_274_5069));
            operation_274_5051 <= ((operation_274_5077)^(operation_274_5070));
            operation_274_5050 <= ((operation_274_5070)^(operation_274_5078));
            operation_274_5049 <= ((operation_274_5069)^(operation_274_5077));
            operation_274_5048 <= ((operation_274_5068)^(operation_274_5074));
            operation_274_5047 <= ((operation_274_5067)^(operation_274_5073));
            operation_274_5046 <= ((operation_274_5066)^(operation_274_5076));
            operation_274_5045 <= ((operation_274_5065)^(operation_274_5075));
            operation_274_5044 <= ((operation_274_5064)^(operation_274_5072));
            operation_274_5043 <= ((operation_274_5063)^(operation_274_5071));
            operation_274_5042 <= ((operation_274_5073)^(operation_274_5068));
            operation_274_5041 <= ((operation_274_5071)^(operation_274_5064));
            operation_274_1536 <= ((operation_274_5164)^(operation_274_1535));
            operation_274_1560 <= ((operation_274_5234)^(operation_274_1655));
            operation_274_5107_latch <= (operation_274_5107);
            operation_274_5106_latch <= (operation_274_5106);
            operation_274_5105_latch <= (operation_274_5105);
            operation_274_5104_latch <= (operation_274_5104);
            operation_274_5103_latch <= (operation_274_5103);
            operation_274_5102_latch <= (operation_274_5102);
            operation_274_5101_latch <= (operation_274_5101);
            operation_274_5100_latch <= (operation_274_5100);
            operation_274_5099_latch <= (operation_274_5099);
            operation_274_5098_latch <= (operation_274_5098);
            operation_274_5097_latch <= (operation_274_5097);
            operation_274_5096_latch <= (operation_274_5096);
            operation_274_5095_latch <= (operation_274_5095);
            operation_274_5094_latch <= (operation_274_5094);
            operation_274_5093_latch <= (operation_274_5093);
            operation_274_5092_latch <= (operation_274_5092);
            operation_274_4304 <= ((operation_274_4322)^(operation_274_4376));
            operation_274_4303 <= ((operation_274_4321)^(operation_274_4375));
            operation_274_4302 <= ((operation_274_4320)^(operation_274_4436));
            operation_274_4301 <= ((operation_274_4319)^(operation_274_4435));
            operation_274_4300 <= ((operation_274_4318)^(operation_274_4496));
            operation_274_4299 <= ((operation_274_4317)^(operation_274_4495));
            operation_274_4298 <= ((operation_274_4316)^(operation_274_4584));
            operation_274_4297 <= ((operation_274_4315)^(operation_274_4583));
            operation_274_4296 <= ((operation_274_4313)^(operation_274_4478));
            operation_274_4295 <= ((operation_274_4312)^(operation_274_4561));
            operation_274_4294 <= ((operation_274_4311)^(operation_274_4418));
            operation_274_4293 <= ((operation_274_4310)^(operation_274_4477));
            operation_274_4292 <= ((operation_274_4309)^(operation_274_4358));
            operation_274_4291 <= ((operation_274_4308)^(operation_274_4417));
            operation_274_4290 <= ((operation_274_4307)^(operation_274_4306));
            operation_274_4289 <= ((operation_274_4305)^(operation_274_4357));
            operation_274_1544 <= ((operation_274_5233)^(operation_274_1639));
            operation_274_1504 <= ((operation_274_5216)^(operation_274_1503));
            operation_274_1552 <= ((operation_274_5215)^(operation_274_1551));
            operation_274_1528 <= ((operation_274_5294)^(operation_274_1623));
            operation_274_4356 <= ((operation_274_4643)^(operation_274_4374));
            operation_274_4355 <= ((operation_274_4642)^(operation_274_4373));
            operation_274_4354 <= ((operation_274_4647)^(operation_274_4372));
            operation_274_4353 <= ((operation_274_4646)^(operation_274_4371));
            operation_274_4352 <= ((operation_274_4645)^(operation_274_4370));
            operation_274_4351 <= ((operation_274_4644)^(operation_274_4369));
            operation_274_4350 <= ((operation_274_4649)^(operation_274_4368));
            operation_274_4349 <= ((operation_274_4648)^(operation_274_4367));
            operation_274_4348 <= ((operation_274_4641)^(operation_274_4366));
            operation_274_4347 <= ((operation_274_4640)^(operation_274_4365));
            operation_274_4346 <= ((operation_274_4639)^(operation_274_4364));
            operation_274_4345 <= ((operation_274_4638)^(operation_274_4363));
            operation_274_4344 <= ((operation_274_4637)^(operation_274_4362));
            operation_274_4343 <= ((operation_274_4636)^(operation_274_4361));
            operation_274_4342 <= ((operation_274_4635)^(operation_274_4360));
            operation_274_4341 <= ((operation_274_4634)^(operation_274_4359));
            operation_274_1512 <= ((operation_274_5293)^(operation_274_1607));
            operation_274_1472 <= ((operation_274_5276)^(operation_274_1471));
            operation_274_1520 <= ((operation_274_5275)^(operation_274_1519));
            operation_274_1496 <= ((operation_274_5354)^(operation_274_1591));
            operation_274_4414 <= ((operation_274_4434)^(operation_274_4499));
            operation_274_4413 <= ((operation_274_4433)^(operation_274_4499));
            operation_274_4412 <= ((operation_274_4432)^(operation_274_4500));
            operation_274_4411 <= ((operation_274_4431)^(operation_274_4500));
            operation_274_4410 <= ((operation_274_4430)^(operation_274_4501));
            operation_274_4409 <= ((operation_274_4429)^(operation_274_4501));
            operation_274_4408 <= ((operation_274_4428)^(operation_274_4502));
            operation_274_4407 <= ((operation_274_4427)^(operation_274_4502));
            operation_274_4406 <= ((operation_274_4426)^(operation_274_4502));
            operation_274_4405 <= ((operation_274_4425)^(operation_274_4502));
            operation_274_4404 <= ((operation_274_4424)^(operation_274_4501));
            operation_274_4403 <= ((operation_274_4423)^(operation_274_4501));
            operation_274_4402 <= ((operation_274_4422)^(operation_274_4500));
            operation_274_4401 <= ((operation_274_4421)^(operation_274_4500));
            operation_274_4400 <= ((operation_274_4420)^(operation_274_4499));
            operation_274_4399 <= ((operation_274_4419)^(operation_274_4499));
            operation_274_1480 <= ((operation_274_5353)^(operation_274_1575));
            operation_274_1440 <= ((operation_274_5336)^(operation_274_1439));
            operation_274_1488 <= ((operation_274_5335)^(operation_274_1487));
            operation_274_1464 <= ((operation_274_5442)^(operation_274_1463));
            operation_274_1423_latch <= (operation_274_1423);
            operation_274_4474 <= ((operation_274_4555)^(operation_274_4494));
            operation_274_4473 <= ((operation_274_4553)^(operation_274_4493));
            operation_274_4472 <= ((operation_274_4551)^(operation_274_4492));
            operation_274_4471 <= ((operation_274_4549)^(operation_274_4491));
            operation_274_4470 <= ((operation_274_4547)^(operation_274_4490));
            operation_274_4469 <= ((operation_274_4545)^(operation_274_4489));
            operation_274_4468 <= ((operation_274_4543)^(operation_274_4488));
            operation_274_4467 <= ((operation_274_4541)^(operation_274_4487));
            operation_274_4466 <= ((operation_274_4540)^(operation_274_4486));
            operation_274_4465 <= ((operation_274_4538)^(operation_274_4485));
            operation_274_4464 <= ((operation_274_4536)^(operation_274_4484));
            operation_274_4463 <= ((operation_274_4534)^(operation_274_4483));
            operation_274_4462 <= ((operation_274_4532)^(operation_274_4482));
            operation_274_4461 <= ((operation_274_4530)^(operation_274_4481));
            operation_274_4460 <= ((operation_274_4528)^(operation_274_4480));
            operation_274_4459 <= ((operation_274_4526)^(operation_274_4479));
            operation_274_1448 <= ((operation_274_5441)^(operation_274_1447));
            operation_274_1432 <= ((operation_274_1428)^(operation_274_5601));
            operation_274_1456 <= ((operation_274_5419)^(operation_274_1455));
            operation_274_4494 <= ((operation_274_4518)*(operation_274_5597));
            operation_274_4493 <= ((operation_274_4517)*(operation_274_5597));
            operation_274_4492 <= ((operation_274_4516)*(operation_274_5597));
            operation_274_4491 <= ((operation_274_4515)*(operation_274_5597));
            operation_274_4490 <= ((operation_274_4514)*(operation_274_5597));
            operation_274_4489 <= ((operation_274_4513)*(operation_274_5597));
            operation_274_4488 <= ((operation_274_4512)*(operation_274_5597));
            operation_274_4487 <= ((operation_274_4511)*(operation_274_5597));
            operation_274_4486 <= ((operation_274_4510)*(operation_274_5597));
            operation_274_4485 <= ((operation_274_4509)*(operation_274_5597));
            operation_274_4484 <= ((operation_274_4508)*(operation_274_5597));
            operation_274_4483 <= ((operation_274_4507)*(operation_274_5597));
            operation_274_4482 <= ((operation_274_4506)*(operation_274_5597));
            operation_274_4481 <= ((operation_274_4505)*(operation_274_5597));
            operation_274_4480 <= ((operation_274_4504)*(operation_274_5597));
            operation_274_4479 <= ((operation_274_4503)*(operation_274_5597));
            operation_274_5198 <= ((operation_274_4735)^(operation_274_5216));
            operation_274_4518 <= ((operation_274_4556)&(operation_274_5557));
            operation_274_4517 <= ((operation_274_4554)&(operation_274_5557));
            operation_274_4516 <= ((operation_274_4552)&(operation_274_5557));
            operation_274_4515 <= ((operation_274_4550)&(operation_274_5557));
            operation_274_4514 <= ((operation_274_4548)&(operation_274_5557));
            operation_274_4513 <= ((operation_274_4546)&(operation_274_5557));
            operation_274_4512 <= ((operation_274_4544)&(operation_274_5557));
            operation_274_4511 <= ((operation_274_4542)&(operation_274_5557));
            operation_274_4510 <= ((operation_274_4539)&(operation_274_5557));
            operation_274_4509 <= ((operation_274_4537)&(operation_274_5557));
            operation_274_4508 <= ((operation_274_4535)&(operation_274_5557));
            operation_274_4507 <= ((operation_274_4533)&(operation_274_5557));
            operation_274_4506 <= ((operation_274_4531)&(operation_274_5557));
            operation_274_4505 <= ((operation_274_4529)&(operation_274_5557));
            operation_274_4504 <= ((operation_274_4527)&(operation_274_5557));
            operation_274_4503 <= ((operation_274_4525)&(operation_274_5557));
            operation_274_1418_latch <= (operation_274_1418);
            operation_274_1408_latch <= (operation_274_1408);
            operation_274_1413_latch <= (operation_274_1413);
            operation_274_4556 <= ((operation_274_4580)>>(operation_274_2119));
            operation_274_4555 <= ((operation_274_4580)<<(operation_274_5557));
            operation_274_4554 <= ((operation_274_4579)>>(operation_274_2119));
            operation_274_4553 <= ((operation_274_4579)<<(operation_274_5557));
            operation_274_4552 <= ((operation_274_4578)>>(operation_274_2119));
            operation_274_4551 <= ((operation_274_4578)<<(operation_274_5557));
            operation_274_4550 <= ((operation_274_4577)>>(operation_274_2119));
            operation_274_4549 <= ((operation_274_4577)<<(operation_274_5557));
            operation_274_4548 <= ((operation_274_4576)>>(operation_274_2119));
            operation_274_4547 <= ((operation_274_4576)<<(operation_274_5557));
            operation_274_4546 <= ((operation_274_4575)>>(operation_274_2119));
            operation_274_4545 <= ((operation_274_4575)<<(operation_274_5557));
            operation_274_4544 <= ((operation_274_4574)>>(operation_274_2119));
            operation_274_4543 <= ((operation_274_4574)<<(operation_274_5557));
            operation_274_4542 <= ((operation_274_4573)>>(operation_274_2119));
            operation_274_4541 <= ((operation_274_4573)<<(operation_274_5557));
            operation_274_4540 <= ((operation_274_4572)<<(operation_274_5557));
            operation_274_4539 <= ((operation_274_4572)>>(operation_274_2119));
            operation_274_4538 <= ((operation_274_4571)<<(operation_274_5557));
            operation_274_4537 <= ((operation_274_4571)>>(operation_274_2119));
            operation_274_4536 <= ((operation_274_4570)<<(operation_274_5557));
            operation_274_4535 <= ((operation_274_4570)>>(operation_274_2119));
            operation_274_4534 <= ((operation_274_4569)<<(operation_274_5557));
            operation_274_4533 <= ((operation_274_4569)>>(operation_274_2119));
            operation_274_4532 <= ((operation_274_4568)<<(operation_274_5557));
            operation_274_4531 <= ((operation_274_4568)>>(operation_274_2119));
            operation_274_4530 <= ((operation_274_4567)<<(operation_274_5557));
            operation_274_4529 <= ((operation_274_4567)>>(operation_274_2119));
            operation_274_4528 <= ((operation_274_4566)<<(operation_274_5557));
            operation_274_4527 <= ((operation_274_4566)>>(operation_274_2119));
            operation_274_4526 <= ((operation_274_4565)<<(operation_274_5557));
            operation_274_4525 <= ((operation_274_4565)>>(operation_274_2119));
            operation_274_4582 <= ((operation_274_4606)^(operation_274_4636));
            operation_274_4581 <= ((operation_274_4605)^(operation_274_4640));
            operation_274_4564 <= ((operation_274_4588)^(operation_274_4638));
            operation_274_4563 <= ((operation_274_4587)^(operation_274_4634));
            operation_274_5274 <= ((operation_274_4805)^(operation_274_5294));
            operation_274_5273 <= ((operation_274_4804)^(operation_274_5293));
            operation_274_5256 <= ((operation_274_4787)^(operation_274_5276));
            operation_274_5255 <= ((operation_274_4786)^(operation_274_5275));
            operation_274_4606 <= ((operation_274_4625)^(operation_274_4647));
            operation_274_4605 <= ((operation_274_4622)^(operation_274_4649));
            operation_274_4588 <= ((operation_274_4613)^(operation_274_4645));
            operation_274_4587 <= ((operation_274_4612)^(operation_274_4643));
            operation_274_4627 <= ((operation_274_4643)^(operation_274_4634));
            operation_274_4626 <= ((operation_274_4647)^(operation_274_4636));
            operation_274_4625 <= ((operation_274_4646)^(operation_274_4637));
            operation_274_4624 <= ((operation_274_4645)^(operation_274_4638));
            operation_274_4623 <= ((operation_274_4649)^(operation_274_4640));
            operation_274_4622 <= ((operation_274_4648)^(operation_274_4641));
            operation_274_4621 <= ((operation_274_4641)^(operation_274_4649));
            operation_274_4620 <= ((operation_274_4640)^(operation_274_4648));
            operation_274_4619 <= ((operation_274_4639)^(operation_274_4645));
            operation_274_4618 <= ((operation_274_4638)^(operation_274_4644));
            operation_274_4617 <= ((operation_274_4637)^(operation_274_4647));
            operation_274_4616 <= ((operation_274_4636)^(operation_274_4646));
            operation_274_4615 <= ((operation_274_4635)^(operation_274_4643));
            operation_274_4614 <= ((operation_274_4634)^(operation_274_4642));
            operation_274_4613 <= ((operation_274_4644)^(operation_274_4639));
            operation_274_4612 <= ((operation_274_4642)^(operation_274_4635));
            operation_274_5334 <= ((operation_274_4865)^(operation_274_5354));
            operation_274_5333 <= ((operation_274_4864)^(operation_274_5353));
            operation_274_5316 <= ((operation_274_4847)^(operation_274_5336));
            operation_274_5315 <= ((operation_274_4846)^(operation_274_5335));
            operation_274_4678_latch <= (operation_274_4678);
            operation_274_4677_latch <= (operation_274_4677);
            operation_274_4676_latch <= (operation_274_4676);
            operation_274_4675_latch <= (operation_274_4675);
            operation_274_4674_latch <= (operation_274_4674);
            operation_274_4673_latch <= (operation_274_4673);
            operation_274_4672_latch <= (operation_274_4672);
            operation_274_4671_latch <= (operation_274_4671);
            operation_274_4670_latch <= (operation_274_4670);
            operation_274_4669_latch <= (operation_274_4669);
            operation_274_4668_latch <= (operation_274_4668);
            operation_274_4667_latch <= (operation_274_4667);
            operation_274_4666_latch <= (operation_274_4666);
            operation_274_4665_latch <= (operation_274_4665);
            operation_274_4664_latch <= (operation_274_4664);
            operation_274_4663_latch <= (operation_274_4663);
            operation_274_3875 <= ((operation_274_3893)^(operation_274_3947));
            operation_274_3874 <= ((operation_274_3892)^(operation_274_3946));
            operation_274_3873 <= ((operation_274_3891)^(operation_274_4007));
            operation_274_3872 <= ((operation_274_3890)^(operation_274_4006));
            operation_274_3871 <= ((operation_274_3889)^(operation_274_4067));
            operation_274_3870 <= ((operation_274_3888)^(operation_274_4066));
            operation_274_3869 <= ((operation_274_3887)^(operation_274_4155));
            operation_274_3868 <= ((operation_274_3886)^(operation_274_4154));
            operation_274_3867 <= ((operation_274_3884)^(operation_274_4049));
            operation_274_3866 <= ((operation_274_3883)^(operation_274_4132));
            operation_274_3865 <= ((operation_274_3882)^(operation_274_3989));
            operation_274_3864 <= ((operation_274_3881)^(operation_274_4048));
            operation_274_3863 <= ((operation_274_3880)^(operation_274_3929));
            operation_274_3862 <= ((operation_274_3879)^(operation_274_3988));
            operation_274_3861 <= ((operation_274_3878)^(operation_274_3877));
            operation_274_3860 <= ((operation_274_3876)^(operation_274_3928));
            operation_274_5418 <= ((operation_274_4925)^(operation_274_5442));
            operation_274_5417 <= ((operation_274_4924)^(operation_274_5441));
            operation_274_5380 <= ((operation_274_4907)^(operation_274_5420));
            operation_274_5379 <= ((operation_274_4906)^(operation_274_5419));
            operation_274_3927 <= ((operation_274_4214)^(operation_274_3945));
            operation_274_3926 <= ((operation_274_4213)^(operation_274_3944));
            operation_274_3925 <= ((operation_274_4218)^(operation_274_3943));
            operation_274_3924 <= ((operation_274_4217)^(operation_274_3942));
            operation_274_3923 <= ((operation_274_4216)^(operation_274_3941));
            operation_274_3922 <= ((operation_274_4215)^(operation_274_3940));
            operation_274_3921 <= ((operation_274_4220)^(operation_274_3939));
            operation_274_3920 <= ((operation_274_4219)^(operation_274_3938));
            operation_274_3919 <= ((operation_274_4212)^(operation_274_3937));
            operation_274_3918 <= ((operation_274_4211)^(operation_274_3936));
            operation_274_3917 <= ((operation_274_4210)^(operation_274_3935));
            operation_274_3916 <= ((operation_274_4209)^(operation_274_3934));
            operation_274_3915 <= ((operation_274_4208)^(operation_274_3933));
            operation_274_3914 <= ((operation_274_4207)^(operation_274_3932));
            operation_274_3913 <= ((operation_274_4206)^(operation_274_3931));
            operation_274_3912 <= ((operation_274_4205)^(operation_274_3930));
            operation_274_5488 <= ((operation_274_5013)^(operation_274_5510));
            operation_274_5487 <= ((operation_274_5012)^(operation_274_5509));
            operation_274_5486 <= ((operation_274_5508)^(operation_274_5597));
            operation_274_5469 <= ((operation_274_4990)^(operation_274_5491));
            operation_274_5538_latch <= (operation_274_5538);
            operation_274_5537_latch <= (operation_274_5537);
            operation_274_5520_latch <= (operation_274_5520);
            operation_274_5519_latch <= (operation_274_5519);
            operation_274_3985 <= ((operation_274_4005)^(operation_274_4070));
            operation_274_3984 <= ((operation_274_4004)^(operation_274_4070));
            operation_274_3983 <= ((operation_274_4003)^(operation_274_4071));
            operation_274_3982 <= ((operation_274_4002)^(operation_274_4071));
            operation_274_3981 <= ((operation_274_4001)^(operation_274_4072));
            operation_274_3980 <= ((operation_274_4000)^(operation_274_4072));
            operation_274_3979 <= ((operation_274_3999)^(operation_274_4073));
            operation_274_3978 <= ((operation_274_3998)^(operation_274_4073));
            operation_274_3977 <= ((operation_274_3997)^(operation_274_4073));
            operation_274_3976 <= ((operation_274_3996)^(operation_274_4073));
            operation_274_3975 <= ((operation_274_3995)^(operation_274_4072));
            operation_274_3974 <= ((operation_274_3994)^(operation_274_4072));
            operation_274_3973 <= ((operation_274_3993)^(operation_274_4071));
            operation_274_3972 <= ((operation_274_3992)^(operation_274_4071));
            operation_274_3971 <= ((operation_274_3991)^(operation_274_4070));
            operation_274_3970 <= ((operation_274_3990)^(operation_274_4070));
            operation_274_4845 <= ((operation_274_4376)^(operation_274_4865));
            operation_274_4844 <= ((operation_274_4375)^(operation_274_4864));
            operation_274_4826 <= ((operation_274_4357)^(operation_274_4846));
            operation_274_4769 <= ((operation_274_4306)^(operation_274_4787));
            operation_274_4045 <= ((operation_274_4126)^(operation_274_4065));
            operation_274_4044 <= ((operation_274_4124)^(operation_274_4064));
            operation_274_4043 <= ((operation_274_4122)^(operation_274_4063));
            operation_274_4042 <= ((operation_274_4120)^(operation_274_4062));
            operation_274_4041 <= ((operation_274_4118)^(operation_274_4061));
            operation_274_4040 <= ((operation_274_4116)^(operation_274_4060));
            operation_274_4039 <= ((operation_274_4114)^(operation_274_4059));
            operation_274_4038 <= ((operation_274_4112)^(operation_274_4058));
            operation_274_4037 <= ((operation_274_4111)^(operation_274_4057));
            operation_274_4036 <= ((operation_274_4109)^(operation_274_4056));
            operation_274_4035 <= ((operation_274_4107)^(operation_274_4055));
            operation_274_4034 <= ((operation_274_4105)^(operation_274_4054));
            operation_274_4033 <= ((operation_274_4103)^(operation_274_4053));
            operation_274_4032 <= ((operation_274_4101)^(operation_274_4052));
            operation_274_4031 <= ((operation_274_4099)^(operation_274_4051));
            operation_274_4030 <= ((operation_274_4097)^(operation_274_4050));
            operation_274_4065 <= ((operation_274_4089)*(operation_274_5597));
            operation_274_4064 <= ((operation_274_4088)*(operation_274_5597));
            operation_274_4063 <= ((operation_274_4087)*(operation_274_5597));
            operation_274_4062 <= ((operation_274_4086)*(operation_274_5597));
            operation_274_4061 <= ((operation_274_4085)*(operation_274_5597));
            operation_274_4060 <= ((operation_274_4084)*(operation_274_5597));
            operation_274_4059 <= ((operation_274_4083)*(operation_274_5597));
            operation_274_4058 <= ((operation_274_4082)*(operation_274_5597));
            operation_274_4057 <= ((operation_274_4081)*(operation_274_5597));
            operation_274_4056 <= ((operation_274_4080)*(operation_274_5597));
            operation_274_4055 <= ((operation_274_4079)*(operation_274_5597));
            operation_274_4054 <= ((operation_274_4078)*(operation_274_5597));
            operation_274_4053 <= ((operation_274_4077)*(operation_274_5597));
            operation_274_4052 <= ((operation_274_4076)*(operation_274_5597));
            operation_274_4051 <= ((operation_274_4075)*(operation_274_5597));
            operation_274_4050 <= ((operation_274_4074)*(operation_274_5597));
            operation_274_4905 <= ((operation_274_4436)^(operation_274_4925));
            operation_274_4904 <= ((operation_274_4435)^(operation_274_4924));
            operation_274_4886 <= ((operation_274_4417)^(operation_274_4906));
            operation_274_4827 <= ((operation_274_4358)^(operation_274_4847));
            operation_274_4089 <= ((operation_274_4127)&(operation_274_5557));
            operation_274_4088 <= ((operation_274_4125)&(operation_274_5557));
            operation_274_4087 <= ((operation_274_4123)&(operation_274_5557));
            operation_274_4086 <= ((operation_274_4121)&(operation_274_5557));
            operation_274_4085 <= ((operation_274_4119)&(operation_274_5557));
            operation_274_4084 <= ((operation_274_4117)&(operation_274_5557));
            operation_274_4083 <= ((operation_274_4115)&(operation_274_5557));
            operation_274_4082 <= ((operation_274_4113)&(operation_274_5557));
            operation_274_4081 <= ((operation_274_4110)&(operation_274_5557));
            operation_274_4080 <= ((operation_274_4108)&(operation_274_5557));
            operation_274_4079 <= ((operation_274_4106)&(operation_274_5557));
            operation_274_4078 <= ((operation_274_4104)&(operation_274_5557));
            operation_274_4077 <= ((operation_274_4102)&(operation_274_5557));
            operation_274_4076 <= ((operation_274_4100)&(operation_274_5557));
            operation_274_4075 <= ((operation_274_4098)&(operation_274_5557));
            operation_274_4074 <= ((operation_274_4096)&(operation_274_5557));
            operation_274_4127 <= ((operation_274_4151)>>(operation_274_2119));
            operation_274_4126 <= ((operation_274_4151)<<(operation_274_5557));
            operation_274_4125 <= ((operation_274_4150)>>(operation_274_2119));
            operation_274_4124 <= ((operation_274_4150)<<(operation_274_5557));
            operation_274_4123 <= ((operation_274_4149)>>(operation_274_2119));
            operation_274_4122 <= ((operation_274_4149)<<(operation_274_5557));
            operation_274_4121 <= ((operation_274_4148)>>(operation_274_2119));
            operation_274_4120 <= ((operation_274_4148)<<(operation_274_5557));
            operation_274_4119 <= ((operation_274_4147)>>(operation_274_2119));
            operation_274_4118 <= ((operation_274_4147)<<(operation_274_5557));
            operation_274_4117 <= ((operation_274_4146)>>(operation_274_2119));
            operation_274_4116 <= ((operation_274_4146)<<(operation_274_5557));
            operation_274_4115 <= ((operation_274_4145)>>(operation_274_2119));
            operation_274_4114 <= ((operation_274_4145)<<(operation_274_5557));
            operation_274_4113 <= ((operation_274_4144)>>(operation_274_2119));
            operation_274_4112 <= ((operation_274_4144)<<(operation_274_5557));
            operation_274_4111 <= ((operation_274_4143)<<(operation_274_5557));
            operation_274_4110 <= ((operation_274_4143)>>(operation_274_2119));
            operation_274_4109 <= ((operation_274_4142)<<(operation_274_5557));
            operation_274_4108 <= ((operation_274_4142)>>(operation_274_2119));
            operation_274_4107 <= ((operation_274_4141)<<(operation_274_5557));
            operation_274_4106 <= ((operation_274_4141)>>(operation_274_2119));
            operation_274_4105 <= ((operation_274_4140)<<(operation_274_5557));
            operation_274_4104 <= ((operation_274_4140)>>(operation_274_2119));
            operation_274_4103 <= ((operation_274_4139)<<(operation_274_5557));
            operation_274_4102 <= ((operation_274_4139)>>(operation_274_2119));
            operation_274_4101 <= ((operation_274_4138)<<(operation_274_5557));
            operation_274_4100 <= ((operation_274_4138)>>(operation_274_2119));
            operation_274_4099 <= ((operation_274_4137)<<(operation_274_5557));
            operation_274_4098 <= ((operation_274_4137)>>(operation_274_2119));
            operation_274_4097 <= ((operation_274_4136)<<(operation_274_5557));
            operation_274_4096 <= ((operation_274_4136)>>(operation_274_2119));
            operation_274_4153 <= ((operation_274_4177)^(operation_274_4207));
            operation_274_4152 <= ((operation_274_4176)^(operation_274_4211));
            operation_274_4135 <= ((operation_274_4159)^(operation_274_4209));
            operation_274_4134 <= ((operation_274_4158)^(operation_274_4205));
            operation_274_4989 <= ((operation_274_4496)^(operation_274_5013));
            operation_274_4988 <= ((operation_274_4495)^(operation_274_5012));
            operation_274_4950 <= ((operation_274_4477)^(operation_274_4990));
            operation_274_4887 <= ((operation_274_4418)^(operation_274_4907));
            operation_274_4177 <= ((operation_274_4196)^(operation_274_4218));
            operation_274_4176 <= ((operation_274_4193)^(operation_274_4220));
            operation_274_4159 <= ((operation_274_4184)^(operation_274_4216));
            operation_274_4158 <= ((operation_274_4183)^(operation_274_4214));
            operation_274_4198 <= ((operation_274_4214)^(operation_274_4205));
            operation_274_4197 <= ((operation_274_4218)^(operation_274_4207));
            operation_274_4196 <= ((operation_274_4217)^(operation_274_4208));
            operation_274_4195 <= ((operation_274_4216)^(operation_274_4209));
            operation_274_4194 <= ((operation_274_4220)^(operation_274_4211));
            operation_274_4193 <= ((operation_274_4219)^(operation_274_4212));
            operation_274_4192 <= ((operation_274_4212)^(operation_274_4220));
            operation_274_4191 <= ((operation_274_4211)^(operation_274_4219));
            operation_274_4190 <= ((operation_274_4210)^(operation_274_4216));
            operation_274_4189 <= ((operation_274_4209)^(operation_274_4215));
            operation_274_4188 <= ((operation_274_4208)^(operation_274_4218));
            operation_274_4187 <= ((operation_274_4207)^(operation_274_4217));
            operation_274_4186 <= ((operation_274_4206)^(operation_274_4214));
            operation_274_4185 <= ((operation_274_4205)^(operation_274_4213));
            operation_274_4184 <= ((operation_274_4215)^(operation_274_4210));
            operation_274_4183 <= ((operation_274_4213)^(operation_274_4206));
            operation_274_5059 <= ((operation_274_4584)^(operation_274_5081));
            operation_274_5058 <= ((operation_274_4583)^(operation_274_5080));
            operation_274_5040 <= ((operation_274_4561)^(operation_274_5062));
            operation_274_4951 <= ((operation_274_4478)^(operation_274_4991));
            operation_274_4249_latch <= (operation_274_4249);
            operation_274_4248_latch <= (operation_274_4248);
            operation_274_4247_latch <= (operation_274_4247);
            operation_274_4246_latch <= (operation_274_4246);
            operation_274_4245_latch <= (operation_274_4245);
            operation_274_4244_latch <= (operation_274_4244);
            operation_274_4243_latch <= (operation_274_4243);
            operation_274_4242_latch <= (operation_274_4242);
            operation_274_4241_latch <= (operation_274_4241);
            operation_274_4240_latch <= (operation_274_4240);
            operation_274_4239_latch <= (operation_274_4239);
            operation_274_4238_latch <= (operation_274_4238);
            operation_274_4237_latch <= (operation_274_4237);
            operation_274_4236_latch <= (operation_274_4236);
            operation_274_4235_latch <= (operation_274_4235);
            operation_274_4234_latch <= (operation_274_4234);
            operation_274_5109_latch <= (operation_274_5109);
            operation_274_5091_latch <= (operation_274_5091);
            operation_274_5090_latch <= (operation_274_5090);
            operation_274_3446 <= ((operation_274_3464)^(operation_274_3518));
            operation_274_3445 <= ((operation_274_3463)^(operation_274_3517));
            operation_274_3444 <= ((operation_274_3462)^(operation_274_3578));
            operation_274_3443 <= ((operation_274_3461)^(operation_274_3577));
            operation_274_3442 <= ((operation_274_3460)^(operation_274_3638));
            operation_274_3441 <= ((operation_274_3459)^(operation_274_3637));
            operation_274_3440 <= ((operation_274_3458)^(operation_274_3726));
            operation_274_3439 <= ((operation_274_3457)^(operation_274_3725));
            operation_274_3438 <= ((operation_274_3455)^(operation_274_3620));
            operation_274_3437 <= ((operation_274_3454)^(operation_274_3703));
            operation_274_3436 <= ((operation_274_3453)^(operation_274_3560));
            operation_274_3435 <= ((operation_274_3452)^(operation_274_3619));
            operation_274_3434 <= ((operation_274_3451)^(operation_274_3500));
            operation_274_3433 <= ((operation_274_3450)^(operation_274_3559));
            operation_274_3432 <= ((operation_274_3449)^(operation_274_3448));
            operation_274_3431 <= ((operation_274_3447)^(operation_274_3499));
            operation_274_5057 <= ((operation_274_5079)^(operation_274_5592));
            operation_274_4416 <= ((operation_274_3947)^(operation_274_4436));
            operation_274_4397 <= ((operation_274_3928)^(operation_274_4417));
            operation_274_4340 <= ((operation_274_3877)^(operation_274_4358));
            operation_274_5108_latch <= (operation_274_5108);
            operation_274_3498 <= ((operation_274_3785)^(operation_274_3516));
            operation_274_3497 <= ((operation_274_3784)^(operation_274_3515));
            operation_274_3496 <= ((operation_274_3789)^(operation_274_3514));
            operation_274_3495 <= ((operation_274_3788)^(operation_274_3513));
            operation_274_3494 <= ((operation_274_3787)^(operation_274_3512));
            operation_274_3493 <= ((operation_274_3786)^(operation_274_3511));
            operation_274_3492 <= ((operation_274_3791)^(operation_274_3510));
            operation_274_3491 <= ((operation_274_3790)^(operation_274_3509));
            operation_274_3490 <= ((operation_274_3783)^(operation_274_3508));
            operation_274_3489 <= ((operation_274_3782)^(operation_274_3507));
            operation_274_3488 <= ((operation_274_3781)^(operation_274_3506));
            operation_274_3487 <= ((operation_274_3780)^(operation_274_3505));
            operation_274_3486 <= ((operation_274_3779)^(operation_274_3504));
            operation_274_3485 <= ((operation_274_3778)^(operation_274_3503));
            operation_274_3484 <= ((operation_274_3777)^(operation_274_3502));
            operation_274_3483 <= ((operation_274_3776)^(operation_274_3501));
            operation_274_4476 <= ((operation_274_4007)^(operation_274_4496));
            operation_274_4457 <= ((operation_274_3988)^(operation_274_4477));
            operation_274_4415 <= ((operation_274_3946)^(operation_274_4435));
            operation_274_4398 <= ((operation_274_3929)^(operation_274_4418));
            operation_274_3556 <= ((operation_274_3576)^(operation_274_3641));
            operation_274_3555 <= ((operation_274_3575)^(operation_274_3641));
            operation_274_3554 <= ((operation_274_3574)^(operation_274_3642));
            operation_274_3553 <= ((operation_274_3573)^(operation_274_3642));
            operation_274_3552 <= ((operation_274_3572)^(operation_274_3643));
            operation_274_3551 <= ((operation_274_3571)^(operation_274_3643));
            operation_274_3550 <= ((operation_274_3570)^(operation_274_3644));
            operation_274_3549 <= ((operation_274_3569)^(operation_274_3644));
            operation_274_3548 <= ((operation_274_3568)^(operation_274_3644));
            operation_274_3547 <= ((operation_274_3567)^(operation_274_3644));
            operation_274_3546 <= ((operation_274_3566)^(operation_274_3643));
            operation_274_3545 <= ((operation_274_3565)^(operation_274_3643));
            operation_274_3544 <= ((operation_274_3564)^(operation_274_3642));
            operation_274_3543 <= ((operation_274_3563)^(operation_274_3642));
            operation_274_3542 <= ((operation_274_3562)^(operation_274_3641));
            operation_274_3541 <= ((operation_274_3561)^(operation_274_3641));
            operation_274_4560 <= ((operation_274_4067)^(operation_274_4584));
            operation_274_4521 <= ((operation_274_4048)^(operation_274_4561));
            operation_274_4475 <= ((operation_274_4006)^(operation_274_4495));
            operation_274_4458 <= ((operation_274_3989)^(operation_274_4478));
            operation_274_3616 <= ((operation_274_3697)^(operation_274_3636));
            operation_274_3615 <= ((operation_274_3695)^(operation_274_3635));
            operation_274_3614 <= ((operation_274_3693)^(operation_274_3634));
            operation_274_3613 <= ((operation_274_3691)^(operation_274_3633));
            operation_274_3612 <= ((operation_274_3689)^(operation_274_3632));
            operation_274_3611 <= ((operation_274_3687)^(operation_274_3631));
            operation_274_3610 <= ((operation_274_3685)^(operation_274_3630));
            operation_274_3609 <= ((operation_274_3683)^(operation_274_3629));
            operation_274_3608 <= ((operation_274_3682)^(operation_274_3628));
            operation_274_3607 <= ((operation_274_3680)^(operation_274_3627));
            operation_274_3606 <= ((operation_274_3678)^(operation_274_3626));
            operation_274_3605 <= ((operation_274_3676)^(operation_274_3625));
            operation_274_3604 <= ((operation_274_3674)^(operation_274_3624));
            operation_274_3603 <= ((operation_274_3672)^(operation_274_3623));
            operation_274_3602 <= ((operation_274_3670)^(operation_274_3622));
            operation_274_3601 <= ((operation_274_3668)^(operation_274_3621));
            operation_274_3636 <= ((operation_274_3660)*(operation_274_5597));
            operation_274_3635 <= ((operation_274_3659)*(operation_274_5597));
            operation_274_3634 <= ((operation_274_3658)*(operation_274_5597));
            operation_274_3633 <= ((operation_274_3657)*(operation_274_5597));
            operation_274_3632 <= ((operation_274_3656)*(operation_274_5597));
            operation_274_3631 <= ((operation_274_3655)*(operation_274_5597));
            operation_274_3630 <= ((operation_274_3654)*(operation_274_5597));
            operation_274_3629 <= ((operation_274_3653)*(operation_274_5597));
            operation_274_3628 <= ((operation_274_3652)*(operation_274_5597));
            operation_274_3627 <= ((operation_274_3651)*(operation_274_5597));
            operation_274_3626 <= ((operation_274_3650)*(operation_274_5597));
            operation_274_3625 <= ((operation_274_3649)*(operation_274_5597));
            operation_274_3624 <= ((operation_274_3648)*(operation_274_5597));
            operation_274_3623 <= ((operation_274_3647)*(operation_274_5597));
            operation_274_3622 <= ((operation_274_3646)*(operation_274_5597));
            operation_274_3621 <= ((operation_274_3645)*(operation_274_5597));
            operation_274_4630 <= ((operation_274_4155)^(operation_274_4652));
            operation_274_4611 <= ((operation_274_4132)^(operation_274_4633));
            operation_274_4559 <= ((operation_274_4066)^(operation_274_4583));
            operation_274_4522 <= ((operation_274_4049)^(operation_274_4562));
            operation_274_3660 <= ((operation_274_3698)&(operation_274_5557));
            operation_274_3659 <= ((operation_274_3696)&(operation_274_5557));
            operation_274_3658 <= ((operation_274_3694)&(operation_274_5557));
            operation_274_3657 <= ((operation_274_3692)&(operation_274_5557));
            operation_274_3656 <= ((operation_274_3690)&(operation_274_5557));
            operation_274_3655 <= ((operation_274_3688)&(operation_274_5557));
            operation_274_3654 <= ((operation_274_3686)&(operation_274_5557));
            operation_274_3653 <= ((operation_274_3684)&(operation_274_5557));
            operation_274_3652 <= ((operation_274_3681)&(operation_274_5557));
            operation_274_3651 <= ((operation_274_3679)&(operation_274_5557));
            operation_274_3650 <= ((operation_274_3677)&(operation_274_5557));
            operation_274_3649 <= ((operation_274_3675)&(operation_274_5557));
            operation_274_3648 <= ((operation_274_3673)&(operation_274_5557));
            operation_274_3647 <= ((operation_274_3671)&(operation_274_5557));
            operation_274_3646 <= ((operation_274_3669)&(operation_274_5557));
            operation_274_3645 <= ((operation_274_3667)&(operation_274_5557));
            operation_274_3698 <= ((operation_274_3722)>>(operation_274_2119));
            operation_274_3697 <= ((operation_274_3722)<<(operation_274_5557));
            operation_274_3696 <= ((operation_274_3721)>>(operation_274_2119));
            operation_274_3695 <= ((operation_274_3721)<<(operation_274_5557));
            operation_274_3694 <= ((operation_274_3720)>>(operation_274_2119));
            operation_274_3693 <= ((operation_274_3720)<<(operation_274_5557));
            operation_274_3692 <= ((operation_274_3719)>>(operation_274_2119));
            operation_274_3691 <= ((operation_274_3719)<<(operation_274_5557));
            operation_274_3690 <= ((operation_274_3718)>>(operation_274_2119));
            operation_274_3689 <= ((operation_274_3718)<<(operation_274_5557));
            operation_274_3688 <= ((operation_274_3717)>>(operation_274_2119));
            operation_274_3687 <= ((operation_274_3717)<<(operation_274_5557));
            operation_274_3686 <= ((operation_274_3716)>>(operation_274_2119));
            operation_274_3685 <= ((operation_274_3716)<<(operation_274_5557));
            operation_274_3684 <= ((operation_274_3715)>>(operation_274_2119));
            operation_274_3683 <= ((operation_274_3715)<<(operation_274_5557));
            operation_274_3682 <= ((operation_274_3714)<<(operation_274_5557));
            operation_274_3681 <= ((operation_274_3714)>>(operation_274_2119));
            operation_274_3680 <= ((operation_274_3713)<<(operation_274_5557));
            operation_274_3679 <= ((operation_274_3713)>>(operation_274_2119));
            operation_274_3678 <= ((operation_274_3712)<<(operation_274_5557));
            operation_274_3677 <= ((operation_274_3712)>>(operation_274_2119));
            operation_274_3676 <= ((operation_274_3711)<<(operation_274_5557));
            operation_274_3675 <= ((operation_274_3711)>>(operation_274_2119));
            operation_274_3674 <= ((operation_274_3710)<<(operation_274_5557));
            operation_274_3673 <= ((operation_274_3710)>>(operation_274_2119));
            operation_274_3672 <= ((operation_274_3709)<<(operation_274_5557));
            operation_274_3671 <= ((operation_274_3709)>>(operation_274_2119));
            operation_274_3670 <= ((operation_274_3708)<<(operation_274_5557));
            operation_274_3669 <= ((operation_274_3708)>>(operation_274_2119));
            operation_274_3668 <= ((operation_274_3707)<<(operation_274_5557));
            operation_274_3667 <= ((operation_274_3707)>>(operation_274_2119));
            operation_274_4680_latch <= (operation_274_4680);
            operation_274_4661_latch <= (operation_274_4661);
            operation_274_3724 <= ((operation_274_3748)^(operation_274_3778));
            operation_274_3723 <= ((operation_274_3747)^(operation_274_3782));
            operation_274_3706 <= ((operation_274_3730)^(operation_274_3780));
            operation_274_3705 <= ((operation_274_3729)^(operation_274_3776));
            operation_274_4629 <= ((operation_274_4154)^(operation_274_4651));
            operation_274_4628 <= ((operation_274_4650)^(operation_274_5587));
            operation_274_3748 <= ((operation_274_3767)^(operation_274_3789));
            operation_274_3747 <= ((operation_274_3764)^(operation_274_3791));
            operation_274_3730 <= ((operation_274_3755)^(operation_274_3787));
            operation_274_3729 <= ((operation_274_3754)^(operation_274_3785));
            operation_274_3987 <= ((operation_274_3518)^(operation_274_4007));
            operation_274_3911 <= ((operation_274_3448)^(operation_274_3929));
            operation_274_3769 <= ((operation_274_3785)^(operation_274_3776));
            operation_274_3768 <= ((operation_274_3789)^(operation_274_3778));
            operation_274_3767 <= ((operation_274_3788)^(operation_274_3779));
            operation_274_3766 <= ((operation_274_3787)^(operation_274_3780));
            operation_274_3765 <= ((operation_274_3791)^(operation_274_3782));
            operation_274_3764 <= ((operation_274_3790)^(operation_274_3783));
            operation_274_3763 <= ((operation_274_3783)^(operation_274_3791));
            operation_274_3762 <= ((operation_274_3782)^(operation_274_3790));
            operation_274_3761 <= ((operation_274_3781)^(operation_274_3787));
            operation_274_3760 <= ((operation_274_3780)^(operation_274_3786));
            operation_274_3759 <= ((operation_274_3779)^(operation_274_3789));
            operation_274_3758 <= ((operation_274_3778)^(operation_274_3788));
            operation_274_3757 <= ((operation_274_3777)^(operation_274_3785));
            operation_274_3756 <= ((operation_274_3776)^(operation_274_3784));
            operation_274_3755 <= ((operation_274_3786)^(operation_274_3781));
            operation_274_3754 <= ((operation_274_3784)^(operation_274_3777));
            operation_274_4679_latch <= (operation_274_4679);
            operation_274_4662_latch <= (operation_274_4662);
            operation_274_3820_latch <= (operation_274_3820);
            operation_274_3819_latch <= (operation_274_3819);
            operation_274_3818_latch <= (operation_274_3818);
            operation_274_3817_latch <= (operation_274_3817);
            operation_274_3816_latch <= (operation_274_3816);
            operation_274_3815_latch <= (operation_274_3815);
            operation_274_3814_latch <= (operation_274_3814);
            operation_274_3813_latch <= (operation_274_3813);
            operation_274_3812_latch <= (operation_274_3812);
            operation_274_3811_latch <= (operation_274_3811);
            operation_274_3810_latch <= (operation_274_3810);
            operation_274_3809_latch <= (operation_274_3809);
            operation_274_3808_latch <= (operation_274_3808);
            operation_274_3807_latch <= (operation_274_3807);
            operation_274_3806_latch <= (operation_274_3806);
            operation_274_3805_latch <= (operation_274_3805);
            operation_274_4047 <= ((operation_274_3578)^(operation_274_4067));
            operation_274_3986 <= ((operation_274_3517)^(operation_274_4006));
            operation_274_3969 <= ((operation_274_3500)^(operation_274_3989));
            operation_274_3968 <= ((operation_274_3499)^(operation_274_3988));
            operation_274_3017 <= ((operation_274_3035)^(operation_274_3089));
            operation_274_3016 <= ((operation_274_3034)^(operation_274_3088));
            operation_274_3015 <= ((operation_274_3033)^(operation_274_3149));
            operation_274_3014 <= ((operation_274_3032)^(operation_274_3148));
            operation_274_3013 <= ((operation_274_3031)^(operation_274_3209));
            operation_274_3012 <= ((operation_274_3030)^(operation_274_3208));
            operation_274_3011 <= ((operation_274_3029)^(operation_274_3297));
            operation_274_3010 <= ((operation_274_3028)^(operation_274_3296));
            operation_274_3009 <= ((operation_274_3026)^(operation_274_3191));
            operation_274_3008 <= ((operation_274_3025)^(operation_274_3274));
            operation_274_3007 <= ((operation_274_3024)^(operation_274_3131));
            operation_274_3006 <= ((operation_274_3023)^(operation_274_3190));
            operation_274_3005 <= ((operation_274_3022)^(operation_274_3071));
            operation_274_3004 <= ((operation_274_3021)^(operation_274_3130));
            operation_274_3003 <= ((operation_274_3020)^(operation_274_3019));
            operation_274_3002 <= ((operation_274_3018)^(operation_274_3070));
            operation_274_4131 <= ((operation_274_3638)^(operation_274_4155));
            operation_274_4046 <= ((operation_274_3577)^(operation_274_4066));
            operation_274_4029 <= ((operation_274_3560)^(operation_274_4049));
            operation_274_4028 <= ((operation_274_3559)^(operation_274_4048));
            operation_274_3069 <= ((operation_274_3356)^(operation_274_3087));
            operation_274_3068 <= ((operation_274_3355)^(operation_274_3086));
            operation_274_3067 <= ((operation_274_3360)^(operation_274_3085));
            operation_274_3066 <= ((operation_274_3359)^(operation_274_3084));
            operation_274_3065 <= ((operation_274_3358)^(operation_274_3083));
            operation_274_3064 <= ((operation_274_3357)^(operation_274_3082));
            operation_274_3063 <= ((operation_274_3362)^(operation_274_3081));
            operation_274_3062 <= ((operation_274_3361)^(operation_274_3080));
            operation_274_3061 <= ((operation_274_3354)^(operation_274_3079));
            operation_274_3060 <= ((operation_274_3353)^(operation_274_3078));
            operation_274_3059 <= ((operation_274_3352)^(operation_274_3077));
            operation_274_3058 <= ((operation_274_3351)^(operation_274_3076));
            operation_274_3057 <= ((operation_274_3350)^(operation_274_3075));
            operation_274_3056 <= ((operation_274_3349)^(operation_274_3074));
            operation_274_3055 <= ((operation_274_3348)^(operation_274_3073));
            operation_274_3054 <= ((operation_274_3347)^(operation_274_3072));
            operation_274_4201 <= ((operation_274_3726)^(operation_274_4223));
            operation_274_4130 <= ((operation_274_3637)^(operation_274_4154));
            operation_274_4093 <= ((operation_274_3620)^(operation_274_4133));
            operation_274_4092 <= ((operation_274_3619)^(operation_274_4132));
            operation_274_3127 <= ((operation_274_3147)^(operation_274_3212));
            operation_274_3126 <= ((operation_274_3146)^(operation_274_3212));
            operation_274_3125 <= ((operation_274_3145)^(operation_274_3213));
            operation_274_3124 <= ((operation_274_3144)^(operation_274_3213));
            operation_274_3123 <= ((operation_274_3143)^(operation_274_3214));
            operation_274_3122 <= ((operation_274_3142)^(operation_274_3214));
            operation_274_3121 <= ((operation_274_3141)^(operation_274_3215));
            operation_274_3120 <= ((operation_274_3140)^(operation_274_3215));
            operation_274_3119 <= ((operation_274_3139)^(operation_274_3215));
            operation_274_3118 <= ((operation_274_3138)^(operation_274_3215));
            operation_274_3117 <= ((operation_274_3137)^(operation_274_3214));
            operation_274_3116 <= ((operation_274_3136)^(operation_274_3214));
            operation_274_3115 <= ((operation_274_3135)^(operation_274_3213));
            operation_274_3114 <= ((operation_274_3134)^(operation_274_3213));
            operation_274_3113 <= ((operation_274_3133)^(operation_274_3212));
            operation_274_3112 <= ((operation_274_3132)^(operation_274_3212));
            operation_274_4232_latch <= (operation_274_4232);
            operation_274_4200 <= ((operation_274_3725)^(operation_274_4222));
            operation_274_4199 <= ((operation_274_4221)^(operation_274_5582));
            operation_274_4182 <= ((operation_274_3703)^(operation_274_4204));
            operation_274_3482 <= ((operation_274_3019)^(operation_274_3500));
            operation_274_3187 <= ((operation_274_3268)^(operation_274_3207));
            operation_274_3186 <= ((operation_274_3266)^(operation_274_3206));
            operation_274_3185 <= ((operation_274_3264)^(operation_274_3205));
            operation_274_3184 <= ((operation_274_3262)^(operation_274_3204));
            operation_274_3183 <= ((operation_274_3260)^(operation_274_3203));
            operation_274_3182 <= ((operation_274_3258)^(operation_274_3202));
            operation_274_3181 <= ((operation_274_3256)^(operation_274_3201));
            operation_274_3180 <= ((operation_274_3254)^(operation_274_3200));
            operation_274_3179 <= ((operation_274_3253)^(operation_274_3199));
            operation_274_3178 <= ((operation_274_3251)^(operation_274_3198));
            operation_274_3177 <= ((operation_274_3249)^(operation_274_3197));
            operation_274_3176 <= ((operation_274_3247)^(operation_274_3196));
            operation_274_3175 <= ((operation_274_3245)^(operation_274_3195));
            operation_274_3174 <= ((operation_274_3243)^(operation_274_3194));
            operation_274_3173 <= ((operation_274_3241)^(operation_274_3193));
            operation_274_3172 <= ((operation_274_3239)^(operation_274_3192));
            operation_274_4251_latch <= (operation_274_4251);
            operation_274_4250_latch <= (operation_274_4250);
            operation_274_4233_latch <= (operation_274_4233);
            operation_274_3207 <= ((operation_274_3231)*(operation_274_5597));
            operation_274_3206 <= ((operation_274_3230)*(operation_274_5597));
            operation_274_3205 <= ((operation_274_3229)*(operation_274_5597));
            operation_274_3204 <= ((operation_274_3228)*(operation_274_5597));
            operation_274_3203 <= ((operation_274_3227)*(operation_274_5597));
            operation_274_3202 <= ((operation_274_3226)*(operation_274_5597));
            operation_274_3201 <= ((operation_274_3225)*(operation_274_5597));
            operation_274_3200 <= ((operation_274_3224)*(operation_274_5597));
            operation_274_3199 <= ((operation_274_3223)*(operation_274_5597));
            operation_274_3198 <= ((operation_274_3222)*(operation_274_5597));
            operation_274_3197 <= ((operation_274_3221)*(operation_274_5597));
            operation_274_3196 <= ((operation_274_3220)*(operation_274_5597));
            operation_274_3195 <= ((operation_274_3219)*(operation_274_5597));
            operation_274_3194 <= ((operation_274_3218)*(operation_274_5597));
            operation_274_3193 <= ((operation_274_3217)*(operation_274_5597));
            operation_274_3192 <= ((operation_274_3216)*(operation_274_5597));
            operation_274_3231 <= ((operation_274_3269)&(operation_274_5557));
            operation_274_3230 <= ((operation_274_3267)&(operation_274_5557));
            operation_274_3229 <= ((operation_274_3265)&(operation_274_5557));
            operation_274_3228 <= ((operation_274_3263)&(operation_274_5557));
            operation_274_3227 <= ((operation_274_3261)&(operation_274_5557));
            operation_274_3226 <= ((operation_274_3259)&(operation_274_5557));
            operation_274_3225 <= ((operation_274_3257)&(operation_274_5557));
            operation_274_3224 <= ((operation_274_3255)&(operation_274_5557));
            operation_274_3223 <= ((operation_274_3252)&(operation_274_5557));
            operation_274_3222 <= ((operation_274_3250)&(operation_274_5557));
            operation_274_3221 <= ((operation_274_3248)&(operation_274_5557));
            operation_274_3220 <= ((operation_274_3246)&(operation_274_5557));
            operation_274_3219 <= ((operation_274_3244)&(operation_274_5557));
            operation_274_3218 <= ((operation_274_3242)&(operation_274_5557));
            operation_274_3217 <= ((operation_274_3240)&(operation_274_5557));
            operation_274_3216 <= ((operation_274_3238)&(operation_274_5557));
            operation_274_3558 <= ((operation_274_3089)^(operation_274_3578));
            operation_274_3557 <= ((operation_274_3088)^(operation_274_3577));
            operation_274_3540 <= ((operation_274_3071)^(operation_274_3560));
            operation_274_3539 <= ((operation_274_3070)^(operation_274_3559));
            operation_274_3269 <= ((operation_274_3293)>>(operation_274_2119));
            operation_274_3268 <= ((operation_274_3293)<<(operation_274_5557));
            operation_274_3267 <= ((operation_274_3292)>>(operation_274_2119));
            operation_274_3266 <= ((operation_274_3292)<<(operation_274_5557));
            operation_274_3265 <= ((operation_274_3291)>>(operation_274_2119));
            operation_274_3264 <= ((operation_274_3291)<<(operation_274_5557));
            operation_274_3263 <= ((operation_274_3290)>>(operation_274_2119));
            operation_274_3262 <= ((operation_274_3290)<<(operation_274_5557));
            operation_274_3261 <= ((operation_274_3289)>>(operation_274_2119));
            operation_274_3260 <= ((operation_274_3289)<<(operation_274_5557));
            operation_274_3259 <= ((operation_274_3288)>>(operation_274_2119));
            operation_274_3258 <= ((operation_274_3288)<<(operation_274_5557));
            operation_274_3257 <= ((operation_274_3287)>>(operation_274_2119));
            operation_274_3256 <= ((operation_274_3287)<<(operation_274_5557));
            operation_274_3255 <= ((operation_274_3286)>>(operation_274_2119));
            operation_274_3254 <= ((operation_274_3286)<<(operation_274_5557));
            operation_274_3253 <= ((operation_274_3285)<<(operation_274_5557));
            operation_274_3252 <= ((operation_274_3285)>>(operation_274_2119));
            operation_274_3251 <= ((operation_274_3284)<<(operation_274_5557));
            operation_274_3250 <= ((operation_274_3284)>>(operation_274_2119));
            operation_274_3249 <= ((operation_274_3283)<<(operation_274_5557));
            operation_274_3248 <= ((operation_274_3283)>>(operation_274_2119));
            operation_274_3247 <= ((operation_274_3282)<<(operation_274_5557));
            operation_274_3246 <= ((operation_274_3282)>>(operation_274_2119));
            operation_274_3245 <= ((operation_274_3281)<<(operation_274_5557));
            operation_274_3244 <= ((operation_274_3281)>>(operation_274_2119));
            operation_274_3243 <= ((operation_274_3280)<<(operation_274_5557));
            operation_274_3242 <= ((operation_274_3280)>>(operation_274_2119));
            operation_274_3241 <= ((operation_274_3279)<<(operation_274_5557));
            operation_274_3240 <= ((operation_274_3279)>>(operation_274_2119));
            operation_274_3239 <= ((operation_274_3278)<<(operation_274_5557));
            operation_274_3238 <= ((operation_274_3278)>>(operation_274_2119));
            operation_274_3295 <= ((operation_274_3319)^(operation_274_3349));
            operation_274_3294 <= ((operation_274_3318)^(operation_274_3353));
            operation_274_3277 <= ((operation_274_3301)^(operation_274_3351));
            operation_274_3276 <= ((operation_274_3300)^(operation_274_3347));
            operation_274_3319 <= ((operation_274_3338)^(operation_274_3360));
            operation_274_3318 <= ((operation_274_3335)^(operation_274_3362));
            operation_274_3301 <= ((operation_274_3326)^(operation_274_3358));
            operation_274_3300 <= ((operation_274_3325)^(operation_274_3356));
            operation_274_3618 <= ((operation_274_3149)^(operation_274_3638));
            operation_274_3617 <= ((operation_274_3148)^(operation_274_3637));
            operation_274_3600 <= ((operation_274_3131)^(operation_274_3620));
            operation_274_3599 <= ((operation_274_3130)^(operation_274_3619));
            operation_274_3340 <= ((operation_274_3356)^(operation_274_3347));
            operation_274_3339 <= ((operation_274_3360)^(operation_274_3349));
            operation_274_3338 <= ((operation_274_3359)^(operation_274_3350));
            operation_274_3337 <= ((operation_274_3358)^(operation_274_3351));
            operation_274_3336 <= ((operation_274_3362)^(operation_274_3353));
            operation_274_3335 <= ((operation_274_3361)^(operation_274_3354));
            operation_274_3334 <= ((operation_274_3354)^(operation_274_3362));
            operation_274_3333 <= ((operation_274_3353)^(operation_274_3361));
            operation_274_3332 <= ((operation_274_3352)^(operation_274_3358));
            operation_274_3331 <= ((operation_274_3351)^(operation_274_3357));
            operation_274_3330 <= ((operation_274_3350)^(operation_274_3360));
            operation_274_3329 <= ((operation_274_3349)^(operation_274_3359));
            operation_274_3328 <= ((operation_274_3348)^(operation_274_3356));
            operation_274_3327 <= ((operation_274_3347)^(operation_274_3355));
            operation_274_3326 <= ((operation_274_3357)^(operation_274_3352));
            operation_274_3325 <= ((operation_274_3355)^(operation_274_3348));
            operation_274_3391_latch <= (operation_274_3391);
            operation_274_3390_latch <= (operation_274_3390);
            operation_274_3389_latch <= (operation_274_3389);
            operation_274_3388_latch <= (operation_274_3388);
            operation_274_3387_latch <= (operation_274_3387);
            operation_274_3386_latch <= (operation_274_3386);
            operation_274_3385_latch <= (operation_274_3385);
            operation_274_3384_latch <= (operation_274_3384);
            operation_274_3383_latch <= (operation_274_3383);
            operation_274_3382_latch <= (operation_274_3382);
            operation_274_3381_latch <= (operation_274_3381);
            operation_274_3380_latch <= (operation_274_3380);
            operation_274_3379_latch <= (operation_274_3379);
            operation_274_3378_latch <= (operation_274_3378);
            operation_274_3377_latch <= (operation_274_3377);
            operation_274_3376_latch <= (operation_274_3376);
            operation_274_3702 <= ((operation_274_3209)^(operation_274_3726));
            operation_274_3701 <= ((operation_274_3208)^(operation_274_3725));
            operation_274_3664 <= ((operation_274_3191)^(operation_274_3704));
            operation_274_3663 <= ((operation_274_3190)^(operation_274_3703));
            operation_274_2588 <= ((operation_274_2606)^(operation_274_2660));
            operation_274_2587 <= ((operation_274_2605)^(operation_274_2659));
            operation_274_2586 <= ((operation_274_2604)^(operation_274_2720));
            operation_274_2585 <= ((operation_274_2603)^(operation_274_2719));
            operation_274_2584 <= ((operation_274_2602)^(operation_274_2780));
            operation_274_2583 <= ((operation_274_2601)^(operation_274_2779));
            operation_274_2582 <= ((operation_274_2600)^(operation_274_2868));
            operation_274_2581 <= ((operation_274_2599)^(operation_274_2867));
            operation_274_2580 <= ((operation_274_2597)^(operation_274_2762));
            operation_274_2579 <= ((operation_274_2596)^(operation_274_2845));
            operation_274_2578 <= ((operation_274_2595)^(operation_274_2702));
            operation_274_2577 <= ((operation_274_2594)^(operation_274_2761));
            operation_274_2576 <= ((operation_274_2593)^(operation_274_2642));
            operation_274_2575 <= ((operation_274_2592)^(operation_274_2701));
            operation_274_2574 <= ((operation_274_2591)^(operation_274_2590));
            operation_274_2573 <= ((operation_274_2589)^(operation_274_2641));
            operation_274_3772 <= ((operation_274_3297)^(operation_274_3794));
            operation_274_3771 <= ((operation_274_3296)^(operation_274_3793));
            operation_274_3770 <= ((operation_274_3792)^(operation_274_5577));
            operation_274_3753 <= ((operation_274_3274)^(operation_274_3775));
            operation_274_2640 <= ((operation_274_2927)^(operation_274_2658));
            operation_274_2639 <= ((operation_274_2926)^(operation_274_2657));
            operation_274_2638 <= ((operation_274_2931)^(operation_274_2656));
            operation_274_2637 <= ((operation_274_2930)^(operation_274_2655));
            operation_274_2636 <= ((operation_274_2929)^(operation_274_2654));
            operation_274_2635 <= ((operation_274_2928)^(operation_274_2653));
            operation_274_2634 <= ((operation_274_2933)^(operation_274_2652));
            operation_274_2633 <= ((operation_274_2932)^(operation_274_2651));
            operation_274_2632 <= ((operation_274_2925)^(operation_274_2650));
            operation_274_2631 <= ((operation_274_2924)^(operation_274_2649));
            operation_274_2630 <= ((operation_274_2923)^(operation_274_2648));
            operation_274_2629 <= ((operation_274_2922)^(operation_274_2647));
            operation_274_2628 <= ((operation_274_2921)^(operation_274_2646));
            operation_274_2627 <= ((operation_274_2920)^(operation_274_2645));
            operation_274_2626 <= ((operation_274_2919)^(operation_274_2644));
            operation_274_2625 <= ((operation_274_2918)^(operation_274_2643));
            operation_274_3822_latch <= (operation_274_3822);
            operation_274_3821_latch <= (operation_274_3821);
            operation_274_3804_latch <= (operation_274_3804);
            operation_274_3803_latch <= (operation_274_3803);
            operation_274_3129 <= ((operation_274_2660)^(operation_274_3149));
            operation_274_3128 <= ((operation_274_2659)^(operation_274_3148));
            operation_274_3110 <= ((operation_274_2641)^(operation_274_3130));
            operation_274_3053 <= ((operation_274_2590)^(operation_274_3071));
            operation_274_2698 <= ((operation_274_2718)^(operation_274_2783));
            operation_274_2697 <= ((operation_274_2717)^(operation_274_2783));
            operation_274_2696 <= ((operation_274_2716)^(operation_274_2784));
            operation_274_2695 <= ((operation_274_2715)^(operation_274_2784));
            operation_274_2694 <= ((operation_274_2714)^(operation_274_2785));
            operation_274_2693 <= ((operation_274_2713)^(operation_274_2785));
            operation_274_2692 <= ((operation_274_2712)^(operation_274_2786));
            operation_274_2691 <= ((operation_274_2711)^(operation_274_2786));
            operation_274_2690 <= ((operation_274_2710)^(operation_274_2786));
            operation_274_2689 <= ((operation_274_2709)^(operation_274_2786));
            operation_274_2688 <= ((operation_274_2708)^(operation_274_2785));
            operation_274_2687 <= ((operation_274_2707)^(operation_274_2785));
            operation_274_2686 <= ((operation_274_2706)^(operation_274_2784));
            operation_274_2685 <= ((operation_274_2705)^(operation_274_2784));
            operation_274_2684 <= ((operation_274_2704)^(operation_274_2783));
            operation_274_2683 <= ((operation_274_2703)^(operation_274_2783));
            operation_274_3189 <= ((operation_274_2720)^(operation_274_3209));
            operation_274_3188 <= ((operation_274_2719)^(operation_274_3208));
            operation_274_3170 <= ((operation_274_2701)^(operation_274_3190));
            operation_274_3111 <= ((operation_274_2642)^(operation_274_3131));
            operation_274_2758 <= ((operation_274_2839)^(operation_274_2778));
            operation_274_2757 <= ((operation_274_2837)^(operation_274_2777));
            operation_274_2756 <= ((operation_274_2835)^(operation_274_2776));
            operation_274_2755 <= ((operation_274_2833)^(operation_274_2775));
            operation_274_2754 <= ((operation_274_2831)^(operation_274_2774));
            operation_274_2753 <= ((operation_274_2829)^(operation_274_2773));
            operation_274_2752 <= ((operation_274_2827)^(operation_274_2772));
            operation_274_2751 <= ((operation_274_2825)^(operation_274_2771));
            operation_274_2750 <= ((operation_274_2824)^(operation_274_2770));
            operation_274_2749 <= ((operation_274_2822)^(operation_274_2769));
            operation_274_2748 <= ((operation_274_2820)^(operation_274_2768));
            operation_274_2747 <= ((operation_274_2818)^(operation_274_2767));
            operation_274_2746 <= ((operation_274_2816)^(operation_274_2766));
            operation_274_2745 <= ((operation_274_2814)^(operation_274_2765));
            operation_274_2744 <= ((operation_274_2812)^(operation_274_2764));
            operation_274_2743 <= ((operation_274_2810)^(operation_274_2763));
            operation_274_2778 <= ((operation_274_2802)*(operation_274_5597));
            operation_274_2777 <= ((operation_274_2801)*(operation_274_5597));
            operation_274_2776 <= ((operation_274_2800)*(operation_274_5597));
            operation_274_2775 <= ((operation_274_2799)*(operation_274_5597));
            operation_274_2774 <= ((operation_274_2798)*(operation_274_5597));
            operation_274_2773 <= ((operation_274_2797)*(operation_274_5597));
            operation_274_2772 <= ((operation_274_2796)*(operation_274_5597));
            operation_274_2771 <= ((operation_274_2795)*(operation_274_5597));
            operation_274_2770 <= ((operation_274_2794)*(operation_274_5597));
            operation_274_2769 <= ((operation_274_2793)*(operation_274_5597));
            operation_274_2768 <= ((operation_274_2792)*(operation_274_5597));
            operation_274_2767 <= ((operation_274_2791)*(operation_274_5597));
            operation_274_2766 <= ((operation_274_2790)*(operation_274_5597));
            operation_274_2765 <= ((operation_274_2789)*(operation_274_5597));
            operation_274_2764 <= ((operation_274_2788)*(operation_274_5597));
            operation_274_2763 <= ((operation_274_2787)*(operation_274_5597));
            operation_274_2802 <= ((operation_274_2840)&(operation_274_5557));
            operation_274_2801 <= ((operation_274_2838)&(operation_274_5557));
            operation_274_2800 <= ((operation_274_2836)&(operation_274_5557));
            operation_274_2799 <= ((operation_274_2834)&(operation_274_5557));
            operation_274_2798 <= ((operation_274_2832)&(operation_274_5557));
            operation_274_2797 <= ((operation_274_2830)&(operation_274_5557));
            operation_274_2796 <= ((operation_274_2828)&(operation_274_5557));
            operation_274_2795 <= ((operation_274_2826)&(operation_274_5557));
            operation_274_2794 <= ((operation_274_2823)&(operation_274_5557));
            operation_274_2793 <= ((operation_274_2821)&(operation_274_5557));
            operation_274_2792 <= ((operation_274_2819)&(operation_274_5557));
            operation_274_2791 <= ((operation_274_2817)&(operation_274_5557));
            operation_274_2790 <= ((operation_274_2815)&(operation_274_5557));
            operation_274_2789 <= ((operation_274_2813)&(operation_274_5557));
            operation_274_2788 <= ((operation_274_2811)&(operation_274_5557));
            operation_274_2787 <= ((operation_274_2809)&(operation_274_5557));
            operation_274_3273 <= ((operation_274_2780)^(operation_274_3297));
            operation_274_3272 <= ((operation_274_2779)^(operation_274_3296));
            operation_274_3234 <= ((operation_274_2761)^(operation_274_3274));
            operation_274_3171 <= ((operation_274_2702)^(operation_274_3191));
            operation_274_2840 <= ((operation_274_2864)>>(operation_274_2119));
            operation_274_2839 <= ((operation_274_2864)<<(operation_274_5557));
            operation_274_2838 <= ((operation_274_2863)>>(operation_274_2119));
            operation_274_2837 <= ((operation_274_2863)<<(operation_274_5557));
            operation_274_2836 <= ((operation_274_2862)>>(operation_274_2119));
            operation_274_2835 <= ((operation_274_2862)<<(operation_274_5557));
            operation_274_2834 <= ((operation_274_2861)>>(operation_274_2119));
            operation_274_2833 <= ((operation_274_2861)<<(operation_274_5557));
            operation_274_2832 <= ((operation_274_2860)>>(operation_274_2119));
            operation_274_2831 <= ((operation_274_2860)<<(operation_274_5557));
            operation_274_2830 <= ((operation_274_2859)>>(operation_274_2119));
            operation_274_2829 <= ((operation_274_2859)<<(operation_274_5557));
            operation_274_2828 <= ((operation_274_2858)>>(operation_274_2119));
            operation_274_2827 <= ((operation_274_2858)<<(operation_274_5557));
            operation_274_2826 <= ((operation_274_2857)>>(operation_274_2119));
            operation_274_2825 <= ((operation_274_2857)<<(operation_274_5557));
            operation_274_2824 <= ((operation_274_2856)<<(operation_274_5557));
            operation_274_2823 <= ((operation_274_2856)>>(operation_274_2119));
            operation_274_2822 <= ((operation_274_2855)<<(operation_274_5557));
            operation_274_2821 <= ((operation_274_2855)>>(operation_274_2119));
            operation_274_2820 <= ((operation_274_2854)<<(operation_274_5557));
            operation_274_2819 <= ((operation_274_2854)>>(operation_274_2119));
            operation_274_2818 <= ((operation_274_2853)<<(operation_274_5557));
            operation_274_2817 <= ((operation_274_2853)>>(operation_274_2119));
            operation_274_2816 <= ((operation_274_2852)<<(operation_274_5557));
            operation_274_2815 <= ((operation_274_2852)>>(operation_274_2119));
            operation_274_2814 <= ((operation_274_2851)<<(operation_274_5557));
            operation_274_2813 <= ((operation_274_2851)>>(operation_274_2119));
            operation_274_2812 <= ((operation_274_2850)<<(operation_274_5557));
            operation_274_2811 <= ((operation_274_2850)>>(operation_274_2119));
            operation_274_2810 <= ((operation_274_2849)<<(operation_274_5557));
            operation_274_2809 <= ((operation_274_2849)>>(operation_274_2119));
            operation_274_2866 <= ((operation_274_2890)^(operation_274_2920));
            operation_274_2865 <= ((operation_274_2889)^(operation_274_2924));
            operation_274_2848 <= ((operation_274_2872)^(operation_274_2922));
            operation_274_2847 <= ((operation_274_2871)^(operation_274_2918));
            operation_274_2890 <= ((operation_274_2909)^(operation_274_2931));
            operation_274_2889 <= ((operation_274_2906)^(operation_274_2933));
            operation_274_2872 <= ((operation_274_2897)^(operation_274_2929));
            operation_274_2871 <= ((operation_274_2896)^(operation_274_2927));
            operation_274_3343 <= ((operation_274_2868)^(operation_274_3365));
            operation_274_3342 <= ((operation_274_2867)^(operation_274_3364));
            operation_274_3324 <= ((operation_274_2845)^(operation_274_3346));
            operation_274_3235 <= ((operation_274_2762)^(operation_274_3275));
            operation_274_2911 <= ((operation_274_2927)^(operation_274_2918));
            operation_274_2910 <= ((operation_274_2931)^(operation_274_2920));
            operation_274_2909 <= ((operation_274_2930)^(operation_274_2921));
            operation_274_2908 <= ((operation_274_2929)^(operation_274_2922));
            operation_274_2907 <= ((operation_274_2933)^(operation_274_2924));
            operation_274_2906 <= ((operation_274_2932)^(operation_274_2925));
            operation_274_2905 <= ((operation_274_2925)^(operation_274_2933));
            operation_274_2904 <= ((operation_274_2924)^(operation_274_2932));
            operation_274_2903 <= ((operation_274_2923)^(operation_274_2929));
            operation_274_2902 <= ((operation_274_2922)^(operation_274_2928));
            operation_274_2901 <= ((operation_274_2921)^(operation_274_2931));
            operation_274_2900 <= ((operation_274_2920)^(operation_274_2930));
            operation_274_2899 <= ((operation_274_2919)^(operation_274_2927));
            operation_274_2898 <= ((operation_274_2918)^(operation_274_2926));
            operation_274_2897 <= ((operation_274_2928)^(operation_274_2923));
            operation_274_2896 <= ((operation_274_2926)^(operation_274_2919));
            operation_274_3393_latch <= (operation_274_3393);
            operation_274_3375_latch <= (operation_274_3375);
            operation_274_3374_latch <= (operation_274_3374);
            operation_274_2962_latch <= (operation_274_2962);
            operation_274_2961_latch <= (operation_274_2961);
            operation_274_2960_latch <= (operation_274_2960);
            operation_274_2959_latch <= (operation_274_2959);
            operation_274_2958_latch <= (operation_274_2958);
            operation_274_2957_latch <= (operation_274_2957);
            operation_274_2956_latch <= (operation_274_2956);
            operation_274_2955_latch <= (operation_274_2955);
            operation_274_2954_latch <= (operation_274_2954);
            operation_274_2953_latch <= (operation_274_2953);
            operation_274_2952_latch <= (operation_274_2952);
            operation_274_2951_latch <= (operation_274_2951);
            operation_274_2950_latch <= (operation_274_2950);
            operation_274_2949_latch <= (operation_274_2949);
            operation_274_2948_latch <= (operation_274_2948);
            operation_274_2947_latch <= (operation_274_2947);
            operation_274_3341 <= ((operation_274_3363)^(operation_274_5572));
            operation_274_2700 <= ((operation_274_2231)^(operation_274_2720));
            operation_274_2681 <= ((operation_274_2212)^(operation_274_2701));
            operation_274_2624 <= ((operation_274_2161)^(operation_274_2642));
            operation_274_2159 <= ((operation_274_2177)^(operation_274_2231));
            operation_274_2158 <= ((operation_274_2176)^(operation_274_2230));
            operation_274_2157 <= ((operation_274_2175)^(operation_274_2291));
            operation_274_2156 <= ((operation_274_2174)^(operation_274_2290));
            operation_274_2155 <= ((operation_274_2173)^(operation_274_2351));
            operation_274_2154 <= ((operation_274_2172)^(operation_274_2350));
            operation_274_2153 <= ((operation_274_2171)^(operation_274_2439));
            operation_274_2152 <= ((operation_274_2170)^(operation_274_2438));
            operation_274_2151 <= ((operation_274_2168)^(operation_274_2333));
            operation_274_2150 <= ((operation_274_2167)^(operation_274_2416));
            operation_274_2149 <= ((operation_274_2166)^(operation_274_2273));
            operation_274_2148 <= ((operation_274_2165)^(operation_274_2332));
            operation_274_2147 <= ((operation_274_2164)^(operation_274_2213));
            operation_274_2146 <= ((operation_274_2163)^(operation_274_2272));
            operation_274_2145 <= ((operation_274_2162)^(operation_274_2161));
            operation_274_2144 <= ((operation_274_2160)^(operation_274_2212));
            operation_274_3392_latch <= (operation_274_3392);
            operation_274_2760 <= ((operation_274_2291)^(operation_274_2780));
            operation_274_2741 <= ((operation_274_2272)^(operation_274_2761));
            operation_274_2699 <= ((operation_274_2230)^(operation_274_2719));
            operation_274_2682 <= ((operation_274_2213)^(operation_274_2702));
            operation_274_2211 <= ((operation_274_2498)^(operation_274_2229));
            operation_274_2210 <= ((operation_274_2497)^(operation_274_2228));
            operation_274_2209 <= ((operation_274_2502)^(operation_274_2227));
            operation_274_2208 <= ((operation_274_2501)^(operation_274_2226));
            operation_274_2207 <= ((operation_274_2500)^(operation_274_2225));
            operation_274_2206 <= ((operation_274_2499)^(operation_274_2224));
            operation_274_2205 <= ((operation_274_2504)^(operation_274_2223));
            operation_274_2204 <= ((operation_274_2503)^(operation_274_2222));
            operation_274_2203 <= ((operation_274_2496)^(operation_274_2221));
            operation_274_2202 <= ((operation_274_2495)^(operation_274_2220));
            operation_274_2201 <= ((operation_274_2494)^(operation_274_2219));
            operation_274_2200 <= ((operation_274_2493)^(operation_274_2218));
            operation_274_2199 <= ((operation_274_2492)^(operation_274_2217));
            operation_274_2198 <= ((operation_274_2491)^(operation_274_2216));
            operation_274_2197 <= ((operation_274_2490)^(operation_274_2215));
            operation_274_2196 <= ((operation_274_2489)^(operation_274_2214));
            operation_274_2844 <= ((operation_274_2351)^(operation_274_2868));
            operation_274_2805 <= ((operation_274_2332)^(operation_274_2845));
            operation_274_2759 <= ((operation_274_2290)^(operation_274_2779));
            operation_274_2742 <= ((operation_274_2273)^(operation_274_2762));
            operation_274_2269 <= ((operation_274_2289)^(operation_274_2354));
            operation_274_2268 <= ((operation_274_2288)^(operation_274_2354));
            operation_274_2267 <= ((operation_274_2287)^(operation_274_2355));
            operation_274_2266 <= ((operation_274_2286)^(operation_274_2355));
            operation_274_2265 <= ((operation_274_2285)^(operation_274_2356));
            operation_274_2264 <= ((operation_274_2284)^(operation_274_2356));
            operation_274_2263 <= ((operation_274_2283)^(operation_274_2357));
            operation_274_2262 <= ((operation_274_2282)^(operation_274_2357));
            operation_274_2261 <= ((operation_274_2281)^(operation_274_2357));
            operation_274_2260 <= ((operation_274_2280)^(operation_274_2357));
            operation_274_2259 <= ((operation_274_2279)^(operation_274_2356));
            operation_274_2258 <= ((operation_274_2278)^(operation_274_2356));
            operation_274_2257 <= ((operation_274_2277)^(operation_274_2355));
            operation_274_2256 <= ((operation_274_2276)^(operation_274_2355));
            operation_274_2255 <= ((operation_274_2275)^(operation_274_2354));
            operation_274_2254 <= ((operation_274_2274)^(operation_274_2354));
            operation_274_2914 <= ((operation_274_2439)^(operation_274_2936));
            operation_274_2895 <= ((operation_274_2416)^(operation_274_2917));
            operation_274_2843 <= ((operation_274_2350)^(operation_274_2867));
            operation_274_2806 <= ((operation_274_2333)^(operation_274_2846));
            operation_274_2329 <= ((operation_274_2410)^(operation_274_2349));
            operation_274_2328 <= ((operation_274_2408)^(operation_274_2348));
            operation_274_2327 <= ((operation_274_2406)^(operation_274_2347));
            operation_274_2326 <= ((operation_274_2404)^(operation_274_2346));
            operation_274_2325 <= ((operation_274_2402)^(operation_274_2345));
            operation_274_2324 <= ((operation_274_2400)^(operation_274_2344));
            operation_274_2323 <= ((operation_274_2398)^(operation_274_2343));
            operation_274_2322 <= ((operation_274_2396)^(operation_274_2342));
            operation_274_2321 <= ((operation_274_2395)^(operation_274_2341));
            operation_274_2320 <= ((operation_274_2393)^(operation_274_2340));
            operation_274_2319 <= ((operation_274_2391)^(operation_274_2339));
            operation_274_2318 <= ((operation_274_2389)^(operation_274_2338));
            operation_274_2317 <= ((operation_274_2387)^(operation_274_2337));
            operation_274_2316 <= ((operation_274_2385)^(operation_274_2336));
            operation_274_2315 <= ((operation_274_2383)^(operation_274_2335));
            operation_274_2314 <= ((operation_274_2381)^(operation_274_2334));
            operation_274_2349 <= ((operation_274_2373)*(operation_274_5597));
            operation_274_2348 <= ((operation_274_2372)*(operation_274_5597));
            operation_274_2347 <= ((operation_274_2371)*(operation_274_5597));
            operation_274_2346 <= ((operation_274_2370)*(operation_274_5597));
            operation_274_2345 <= ((operation_274_2369)*(operation_274_5597));
            operation_274_2344 <= ((operation_274_2368)*(operation_274_5597));
            operation_274_2343 <= ((operation_274_2367)*(operation_274_5597));
            operation_274_2342 <= ((operation_274_2366)*(operation_274_5597));
            operation_274_2341 <= ((operation_274_2365)*(operation_274_5597));
            operation_274_2340 <= ((operation_274_2364)*(operation_274_5597));
            operation_274_2339 <= ((operation_274_2363)*(operation_274_5597));
            operation_274_2338 <= ((operation_274_2362)*(operation_274_5597));
            operation_274_2337 <= ((operation_274_2361)*(operation_274_5597));
            operation_274_2336 <= ((operation_274_2360)*(operation_274_5597));
            operation_274_2335 <= ((operation_274_2359)*(operation_274_5597));
            operation_274_2334 <= ((operation_274_2358)*(operation_274_5597));
            operation_274_2964_latch <= (operation_274_2964);
            operation_274_2945_latch <= (operation_274_2945);
            operation_274_2373 <= ((operation_274_2411)&(operation_274_5557));
            operation_274_2372 <= ((operation_274_2409)&(operation_274_5557));
            operation_274_2371 <= ((operation_274_2407)&(operation_274_5557));
            operation_274_2370 <= ((operation_274_2405)&(operation_274_5557));
            operation_274_2369 <= ((operation_274_2403)&(operation_274_5557));
            operation_274_2368 <= ((operation_274_2401)&(operation_274_5557));
            operation_274_2367 <= ((operation_274_2399)&(operation_274_5557));
            operation_274_2366 <= ((operation_274_2397)&(operation_274_5557));
            operation_274_2365 <= ((operation_274_2394)&(operation_274_5557));
            operation_274_2364 <= ((operation_274_2392)&(operation_274_5557));
            operation_274_2363 <= ((operation_274_2390)&(operation_274_5557));
            operation_274_2362 <= ((operation_274_2388)&(operation_274_5557));
            operation_274_2361 <= ((operation_274_2386)&(operation_274_5557));
            operation_274_2360 <= ((operation_274_2384)&(operation_274_5557));
            operation_274_2359 <= ((operation_274_2382)&(operation_274_5557));
            operation_274_2358 <= ((operation_274_2380)&(operation_274_5557));
            operation_274_2913 <= ((operation_274_2438)^(operation_274_2935));
            operation_274_2912 <= ((operation_274_2934)^(operation_274_5567));
            operation_274_2411 <= ((operation_274_2435)>>(operation_274_2119));
            operation_274_2410 <= ((operation_274_2435)<<(operation_274_5557));
            operation_274_2409 <= ((operation_274_2434)>>(operation_274_2119));
            operation_274_2408 <= ((operation_274_2434)<<(operation_274_5557));
            operation_274_2407 <= ((operation_274_2433)>>(operation_274_2119));
            operation_274_2406 <= ((operation_274_2433)<<(operation_274_5557));
            operation_274_2405 <= ((operation_274_2432)>>(operation_274_2119));
            operation_274_2404 <= ((operation_274_2432)<<(operation_274_5557));
            operation_274_2403 <= ((operation_274_2431)>>(operation_274_2119));
            operation_274_2402 <= ((operation_274_2431)<<(operation_274_5557));
            operation_274_2401 <= ((operation_274_2430)>>(operation_274_2119));
            operation_274_2400 <= ((operation_274_2430)<<(operation_274_5557));
            operation_274_2399 <= ((operation_274_2429)>>(operation_274_2119));
            operation_274_2398 <= ((operation_274_2429)<<(operation_274_5557));
            operation_274_2397 <= ((operation_274_2428)>>(operation_274_2119));
            operation_274_2396 <= ((operation_274_2428)<<(operation_274_5557));
            operation_274_2395 <= ((operation_274_2427)<<(operation_274_5557));
            operation_274_2394 <= ((operation_274_2427)>>(operation_274_2119));
            operation_274_2393 <= ((operation_274_2426)<<(operation_274_5557));
            operation_274_2392 <= ((operation_274_2426)>>(operation_274_2119));
            operation_274_2391 <= ((operation_274_2425)<<(operation_274_5557));
            operation_274_2390 <= ((operation_274_2425)>>(operation_274_2119));
            operation_274_2389 <= ((operation_274_2424)<<(operation_274_5557));
            operation_274_2388 <= ((operation_274_2424)>>(operation_274_2119));
            operation_274_2387 <= ((operation_274_2423)<<(operation_274_5557));
            operation_274_2386 <= ((operation_274_2423)>>(operation_274_2119));
            operation_274_2385 <= ((operation_274_2422)<<(operation_274_5557));
            operation_274_2384 <= ((operation_274_2422)>>(operation_274_2119));
            operation_274_2383 <= ((operation_274_2421)<<(operation_274_5557));
            operation_274_2382 <= ((operation_274_2421)>>(operation_274_2119));
            operation_274_2381 <= ((operation_274_2420)<<(operation_274_5557));
            operation_274_2380 <= ((operation_274_2420)>>(operation_274_2119));
            operation_274_2271 <= ((operation_274_1802)^(operation_274_2291));
            operation_274_2195 <= ((operation_274_1732)^(operation_274_2213));
            operation_274_2437 <= ((operation_274_2461)^(operation_274_2491));
            operation_274_2436 <= ((operation_274_2460)^(operation_274_2495));
            operation_274_2419 <= ((operation_274_2443)^(operation_274_2493));
            operation_274_2418 <= ((operation_274_2442)^(operation_274_2489));
            operation_274_2963_latch <= (operation_274_2963);
            operation_274_2946_latch <= (operation_274_2946);
            operation_274_2461 <= ((operation_274_2480)^(operation_274_2502));
            operation_274_2460 <= ((operation_274_2477)^(operation_274_2504));
            operation_274_2443 <= ((operation_274_2468)^(operation_274_2500));
            operation_274_2442 <= ((operation_274_2467)^(operation_274_2498));
            operation_274_2482 <= ((operation_274_2498)^(operation_274_2489));
            operation_274_2481 <= ((operation_274_2502)^(operation_274_2491));
            operation_274_2480 <= ((operation_274_2501)^(operation_274_2492));
            operation_274_2479 <= ((operation_274_2500)^(operation_274_2493));
            operation_274_2478 <= ((operation_274_2504)^(operation_274_2495));
            operation_274_2477 <= ((operation_274_2503)^(operation_274_2496));
            operation_274_2476 <= ((operation_274_2496)^(operation_274_2504));
            operation_274_2475 <= ((operation_274_2495)^(operation_274_2503));
            operation_274_2474 <= ((operation_274_2494)^(operation_274_2500));
            operation_274_2473 <= ((operation_274_2493)^(operation_274_2499));
            operation_274_2472 <= ((operation_274_2492)^(operation_274_2502));
            operation_274_2471 <= ((operation_274_2491)^(operation_274_2501));
            operation_274_2470 <= ((operation_274_2490)^(operation_274_2498));
            operation_274_2469 <= ((operation_274_2489)^(operation_274_2497));
            operation_274_2468 <= ((operation_274_2499)^(operation_274_2494));
            operation_274_2467 <= ((operation_274_2497)^(operation_274_2490));
            operation_274_2331 <= ((operation_274_1862)^(operation_274_2351));
            operation_274_2270 <= ((operation_274_1801)^(operation_274_2290));
            operation_274_2253 <= ((operation_274_1784)^(operation_274_2273));
            operation_274_2252 <= ((operation_274_1783)^(operation_274_2272));
            operation_274_2533_latch <= (operation_274_2533);
            operation_274_2532_latch <= (operation_274_2532);
            operation_274_2531_latch <= (operation_274_2531);
            operation_274_2530_latch <= (operation_274_2530);
            operation_274_2529_latch <= (operation_274_2529);
            operation_274_2528_latch <= (operation_274_2528);
            operation_274_2527_latch <= (operation_274_2527);
            operation_274_2526_latch <= (operation_274_2526);
            operation_274_2525_latch <= (operation_274_2525);
            operation_274_2524_latch <= (operation_274_2524);
            operation_274_2523_latch <= (operation_274_2523);
            operation_274_2522_latch <= (operation_274_2522);
            operation_274_2521_latch <= (operation_274_2521);
            operation_274_2520_latch <= (operation_274_2520);
            operation_274_2519_latch <= (operation_274_2519);
            operation_274_2518_latch <= (operation_274_2518);
            operation_274_2415 <= ((operation_274_1922)^(operation_274_2439));
            operation_274_2330 <= ((operation_274_1861)^(operation_274_2350));
            operation_274_2313 <= ((operation_274_1844)^(operation_274_2333));
            operation_274_2312 <= ((operation_274_1843)^(operation_274_2332));
            operation_274_1730 <= ((operation_274_1748)^(operation_274_1802));
            operation_274_1729 <= ((operation_274_1747)^(operation_274_1801));
            operation_274_1728 <= ((operation_274_1746)^(operation_274_1862));
            operation_274_1727 <= ((operation_274_1745)^(operation_274_1861));
            operation_274_1726 <= ((operation_274_1744)^(operation_274_1922));
            operation_274_1725 <= ((operation_274_1743)^(operation_274_1921));
            operation_274_1724 <= ((operation_274_1742)^(operation_274_2010));
            operation_274_1723 <= ((operation_274_1741)^(operation_274_2009));
            operation_274_1722 <= ((operation_274_1739)^(operation_274_1904));
            operation_274_1721 <= ((operation_274_1738)^(operation_274_1987));
            operation_274_1720 <= ((operation_274_1737)^(operation_274_1844));
            operation_274_1719 <= ((operation_274_1736)^(operation_274_1903));
            operation_274_1718 <= ((operation_274_1735)^(operation_274_1784));
            operation_274_1717 <= ((operation_274_1734)^(operation_274_1843));
            operation_274_1716 <= ((operation_274_1733)^(operation_274_1732));
            operation_274_1715 <= ((operation_274_1731)^(operation_274_1783));
            operation_274_2485 <= ((operation_274_2010)^(operation_274_2507));
            operation_274_2414 <= ((operation_274_1921)^(operation_274_2438));
            operation_274_2377 <= ((operation_274_1904)^(operation_274_2417));
            operation_274_2376 <= ((operation_274_1903)^(operation_274_2416));
            operation_274_1782 <= ((operation_274_2069)^(operation_274_1800));
            operation_274_1781 <= ((operation_274_2068)^(operation_274_1799));
            operation_274_1780 <= ((operation_274_2073)^(operation_274_1798));
            operation_274_1779 <= ((operation_274_2072)^(operation_274_1797));
            operation_274_1778 <= ((operation_274_2071)^(operation_274_1796));
            operation_274_1777 <= ((operation_274_2070)^(operation_274_1795));
            operation_274_1776 <= ((operation_274_2075)^(operation_274_1794));
            operation_274_1775 <= ((operation_274_2074)^(operation_274_1793));
            operation_274_1774 <= ((operation_274_2067)^(operation_274_1792));
            operation_274_1773 <= ((operation_274_2066)^(operation_274_1791));
            operation_274_1772 <= ((operation_274_2065)^(operation_274_1790));
            operation_274_1771 <= ((operation_274_2064)^(operation_274_1789));
            operation_274_1770 <= ((operation_274_2063)^(operation_274_1788));
            operation_274_1769 <= ((operation_274_2062)^(operation_274_1787));
            operation_274_1768 <= ((operation_274_2061)^(operation_274_1786));
            operation_274_1767 <= ((operation_274_2060)^(operation_274_1785));
            operation_274_2516_latch <= (operation_274_2516);
            operation_274_2484 <= ((operation_274_2009)^(operation_274_2506));
            operation_274_2483 <= ((operation_274_2505)^(operation_274_5562));
            operation_274_2466 <= ((operation_274_1987)^(operation_274_2488));
            operation_274_1840 <= ((operation_274_1860)^(operation_274_1925));
            operation_274_1839 <= ((operation_274_1859)^(operation_274_1925));
            operation_274_1838 <= ((operation_274_1858)^(operation_274_1926));
            operation_274_1837 <= ((operation_274_1857)^(operation_274_1926));
            operation_274_1836 <= ((operation_274_1856)^(operation_274_1927));
            operation_274_1835 <= ((operation_274_1855)^(operation_274_1927));
            operation_274_1834 <= ((operation_274_1854)^(operation_274_1928));
            operation_274_1833 <= ((operation_274_1853)^(operation_274_1928));
            operation_274_1832 <= ((operation_274_1852)^(operation_274_1928));
            operation_274_1831 <= ((operation_274_1851)^(operation_274_1928));
            operation_274_1830 <= ((operation_274_1850)^(operation_274_1927));
            operation_274_1829 <= ((operation_274_1849)^(operation_274_1927));
            operation_274_1828 <= ((operation_274_1848)^(operation_274_1926));
            operation_274_1827 <= ((operation_274_1847)^(operation_274_1926));
            operation_274_1826 <= ((operation_274_1846)^(operation_274_1925));
            operation_274_1825 <= ((operation_274_1845)^(operation_274_1925));
            operation_274_1766 <= ((operation_274_101)^(operation_274_1784));
            operation_274_2535_latch <= (operation_274_2535);
            operation_274_2534_latch <= (operation_274_2534);
            operation_274_2517_latch <= (operation_274_2517);
            operation_274_1900 <= ((operation_274_1981)^(operation_274_1920));
            operation_274_1899 <= ((operation_274_1979)^(operation_274_1919));
            operation_274_1898 <= ((operation_274_1977)^(operation_274_1918));
            operation_274_1897 <= ((operation_274_1975)^(operation_274_1917));
            operation_274_1896 <= ((operation_274_1973)^(operation_274_1916));
            operation_274_1895 <= ((operation_274_1971)^(operation_274_1915));
            operation_274_1894 <= ((operation_274_1969)^(operation_274_1914));
            operation_274_1893 <= ((operation_274_1967)^(operation_274_1913));
            operation_274_1892 <= ((operation_274_1966)^(operation_274_1912));
            operation_274_1891 <= ((operation_274_1964)^(operation_274_1911));
            operation_274_1890 <= ((operation_274_1962)^(operation_274_1910));
            operation_274_1889 <= ((operation_274_1960)^(operation_274_1909));
            operation_274_1888 <= ((operation_274_1958)^(operation_274_1908));
            operation_274_1887 <= ((operation_274_1956)^(operation_274_1907));
            operation_274_1886 <= ((operation_274_1954)^(operation_274_1906));
            operation_274_1885 <= ((operation_274_1952)^(operation_274_1905));
            operation_274_1842 <= ((operation_274_125)^(operation_274_1862));
            operation_274_1841 <= ((operation_274_109)^(operation_274_1861));
            operation_274_1824 <= ((operation_274_69)^(operation_274_1844));
            operation_274_1823 <= ((operation_274_117)^(operation_274_1843));
            operation_274_1920 <= ((operation_274_1944)*(operation_274_5597));
            operation_274_1919 <= ((operation_274_1943)*(operation_274_5597));
            operation_274_1918 <= ((operation_274_1942)*(operation_274_5597));
            operation_274_1917 <= ((operation_274_1941)*(operation_274_5597));
            operation_274_1916 <= ((operation_274_1940)*(operation_274_5597));
            operation_274_1915 <= ((operation_274_1939)*(operation_274_5597));
            operation_274_1914 <= ((operation_274_1938)*(operation_274_5597));
            operation_274_1913 <= ((operation_274_1937)*(operation_274_5597));
            operation_274_1912 <= ((operation_274_1936)*(operation_274_5597));
            operation_274_1911 <= ((operation_274_1935)*(operation_274_5597));
            operation_274_1910 <= ((operation_274_1934)*(operation_274_5597));
            operation_274_1909 <= ((operation_274_1933)*(operation_274_5597));
            operation_274_1908 <= ((operation_274_1932)*(operation_274_5597));
            operation_274_1907 <= ((operation_274_1931)*(operation_274_5597));
            operation_274_1906 <= ((operation_274_1930)*(operation_274_5597));
            operation_274_1905 <= ((operation_274_1929)*(operation_274_5597));
            operation_274_1944 <= ((operation_274_1982)&(operation_274_5557));
            operation_274_1943 <= ((operation_274_1980)&(operation_274_5557));
            operation_274_1942 <= ((operation_274_1978)&(operation_274_5557));
            operation_274_1941 <= ((operation_274_1976)&(operation_274_5557));
            operation_274_1940 <= ((operation_274_1974)&(operation_274_5557));
            operation_274_1939 <= ((operation_274_1972)&(operation_274_5557));
            operation_274_1938 <= ((operation_274_1970)&(operation_274_5557));
            operation_274_1937 <= ((operation_274_1968)&(operation_274_5557));
            operation_274_1936 <= ((operation_274_1965)&(operation_274_5557));
            operation_274_1935 <= ((operation_274_1963)&(operation_274_5557));
            operation_274_1934 <= ((operation_274_1961)&(operation_274_5557));
            operation_274_1933 <= ((operation_274_1959)&(operation_274_5557));
            operation_274_1932 <= ((operation_274_1957)&(operation_274_5557));
            operation_274_1931 <= ((operation_274_1955)&(operation_274_5557));
            operation_274_1930 <= ((operation_274_1953)&(operation_274_5557));
            operation_274_1929 <= ((operation_274_1951)&(operation_274_5557));
            operation_274_1982 <= ((operation_274_2006)>>(operation_274_2119));
            operation_274_1981 <= ((operation_274_2006)<<(operation_274_5557));
            operation_274_1980 <= ((operation_274_2005)>>(operation_274_2119));
            operation_274_1979 <= ((operation_274_2005)<<(operation_274_5557));
            operation_274_1978 <= ((operation_274_2004)>>(operation_274_2119));
            operation_274_1977 <= ((operation_274_2004)<<(operation_274_5557));
            operation_274_1976 <= ((operation_274_2003)>>(operation_274_2119));
            operation_274_1975 <= ((operation_274_2003)<<(operation_274_5557));
            operation_274_1974 <= ((operation_274_2002)>>(operation_274_2119));
            operation_274_1973 <= ((operation_274_2002)<<(operation_274_5557));
            operation_274_1972 <= ((operation_274_2001)>>(operation_274_2119));
            operation_274_1971 <= ((operation_274_2001)<<(operation_274_5557));
            operation_274_1970 <= ((operation_274_2000)>>(operation_274_2119));
            operation_274_1969 <= ((operation_274_2000)<<(operation_274_5557));
            operation_274_1968 <= ((operation_274_1999)>>(operation_274_2119));
            operation_274_1967 <= ((operation_274_1999)<<(operation_274_5557));
            operation_274_1966 <= ((operation_274_1998)<<(operation_274_5557));
            operation_274_1965 <= ((operation_274_1998)>>(operation_274_2119));
            operation_274_1964 <= ((operation_274_1997)<<(operation_274_5557));
            operation_274_1963 <= ((operation_274_1997)>>(operation_274_2119));
            operation_274_1962 <= ((operation_274_1996)<<(operation_274_5557));
            operation_274_1961 <= ((operation_274_1996)>>(operation_274_2119));
            operation_274_1960 <= ((operation_274_1995)<<(operation_274_5557));
            operation_274_1959 <= ((operation_274_1995)>>(operation_274_2119));
            operation_274_1958 <= ((operation_274_1994)<<(operation_274_5557));
            operation_274_1957 <= ((operation_274_1994)>>(operation_274_2119));
            operation_274_1956 <= ((operation_274_1993)<<(operation_274_5557));
            operation_274_1955 <= ((operation_274_1993)>>(operation_274_2119));
            operation_274_1954 <= ((operation_274_1992)<<(operation_274_5557));
            operation_274_1953 <= ((operation_274_1992)>>(operation_274_2119));
            operation_274_1952 <= ((operation_274_1991)<<(operation_274_5557));
            operation_274_1951 <= ((operation_274_1991)>>(operation_274_2119));
            operation_274_1902 <= ((operation_274_93)^(operation_274_1922));
            operation_274_1901 <= ((operation_274_77)^(operation_274_1921));
            operation_274_1884 <= ((operation_274_37)^(operation_274_1904));
            operation_274_1883 <= ((operation_274_85)^(operation_274_1903));
            operation_274_2008 <= ((operation_274_2032)^(operation_274_2062));
            operation_274_2007 <= ((operation_274_2031)^(operation_274_2066));
            operation_274_1990 <= ((operation_274_2014)^(operation_274_2064));
            operation_274_1989 <= ((operation_274_2013)^(operation_274_2060));
            operation_274_2032 <= ((operation_274_2051)^(operation_274_2073));
            operation_274_2031 <= ((operation_274_2048)^(operation_274_2075));
            operation_274_2014 <= ((operation_274_2039)^(operation_274_2071));
            operation_274_2013 <= ((operation_274_2038)^(operation_274_2069));
            operation_274_2053 <= ((operation_274_2069)^(operation_274_2060));
            operation_274_2052 <= ((operation_274_2073)^(operation_274_2062));
            operation_274_2051 <= ((operation_274_2072)^(operation_274_2063));
            operation_274_2050 <= ((operation_274_2071)^(operation_274_2064));
            operation_274_2049 <= ((operation_274_2075)^(operation_274_2066));
            operation_274_2048 <= ((operation_274_2074)^(operation_274_2067));
            operation_274_2047 <= ((operation_274_2067)^(operation_274_2075));
            operation_274_2046 <= ((operation_274_2066)^(operation_274_2074));
            operation_274_2045 <= ((operation_274_2065)^(operation_274_2071));
            operation_274_2044 <= ((operation_274_2064)^(operation_274_2070));
            operation_274_2043 <= ((operation_274_2063)^(operation_274_2073));
            operation_274_2042 <= ((operation_274_2062)^(operation_274_2072));
            operation_274_2041 <= ((operation_274_2061)^(operation_274_2069));
            operation_274_2040 <= ((operation_274_2060)^(operation_274_2068));
            operation_274_2039 <= ((operation_274_2070)^(operation_274_2065));
            operation_274_2038 <= ((operation_274_2068)^(operation_274_2061));
            operation_274_1986 <= ((operation_274_61)^(operation_274_2010));
            operation_274_1985 <= ((operation_274_45)^(operation_274_2009));
            operation_274_1948 <= ((operation_274_5)^(operation_274_1988));
            operation_274_1947 <= ((operation_274_53)^(operation_274_1987));
            operation_274_2104_latch <= (operation_274_2104);
            operation_274_2103_latch <= (operation_274_2103);
            operation_274_2102_latch <= (operation_274_2102);
            operation_274_2101_latch <= (operation_274_2101);
            operation_274_2100_latch <= (operation_274_2100);
            operation_274_2099_latch <= (operation_274_2099);
            operation_274_2098_latch <= (operation_274_2098);
            operation_274_2097_latch <= (operation_274_2097);
            operation_274_2096_latch <= (operation_274_2096);
            operation_274_2095_latch <= (operation_274_2095);
            operation_274_2094_latch <= (operation_274_2094);
            operation_274_2093_latch <= (operation_274_2093);
            operation_274_2092_latch <= (operation_274_2092);
            operation_274_2091_latch <= (operation_274_2091);
            operation_274_2090_latch <= (operation_274_2090);
            operation_274_2089_latch <= (operation_274_2089);
            operation_274_2056 <= ((operation_274_29)^(operation_274_2078));
            operation_274_2055 <= ((operation_274_13)^(operation_274_2077));
            operation_274_2054 <= ((operation_274_2076)^(operation_274_5557));
            operation_274_2037 <= ((operation_274_21)^(operation_274_2059));
            operation_274_118 <= ((operation_274_115)^(operation_274_117));
            operation_274_102 <= ((operation_274_99)^(operation_274_101));
            operation_274_86 <= ((operation_274_83)^(operation_274_85));
            operation_274_70 <= ((operation_274_67)^(operation_274_69));
            operation_274_54 <= ((operation_274_51)^(operation_274_53));
            operation_274_38 <= ((operation_274_35)^(operation_274_37));
            operation_274_22 <= ((operation_274_19)^(operation_274_21));
            operation_274_6 <= ((operation_274_3)^(operation_274_5));
            operation_274_14 <= ((operation_274_11)^(operation_274_13));
            operation_274_30 <= ((operation_274_27)^(operation_274_29));
            operation_274_46 <= ((operation_274_43)^(operation_274_45));
            operation_274_62 <= ((operation_274_59)^(operation_274_61));
            operation_274_78 <= ((operation_274_75)^(operation_274_77));
            operation_274_94 <= ((operation_274_91)^(operation_274_93));
            operation_274_110 <= ((operation_274_107)^(operation_274_109));
            operation_274_126 <= ((operation_274_123)^(operation_274_125));
            operation_274_2106_latch <= (operation_274_2106);
            operation_274_2105_latch <= (operation_274_2105);
            operation_274_2088_latch <= (operation_274_2088);
            operation_274_2087_latch <= (operation_274_2087);
            control_274_follow <= (control_274_end);
            control_274_84 <= (control_274_83);
            control_274_83 <= (control_274_82);
            control_274_82 <= (control_274_81);
            control_274_81 <= (control_274_80);
            control_274_80 <= (control_274_79);
            control_274_79 <= (control_274_78);
            control_274_78 <= (control_274_77);
            control_274_77 <= (control_274_76);
            control_274_76 <= (control_274_75);
            control_274_75 <= (control_274_74);
            control_274_74 <= (control_274_73);
            control_274_73 <= (control_274_72);
            control_274_72 <= (control_274_71);
            control_274_71 <= (control_274_70);
            control_274_70 <= (control_274_69);
            control_274_69 <= (control_274_68);
            control_274_68 <= (control_274_67);
            control_274_67 <= (control_274_66);
            control_274_66 <= (control_274_65);
            control_274_65 <= (control_274_64);
            control_274_64 <= (control_274_63);
            control_274_63 <= (control_274_62);
            control_274_62 <= (control_274_61);
            control_274_61 <= (control_274_60);
            control_274_60 <= (control_274_59);
            control_274_59 <= (control_274_58);
            control_274_58 <= (control_274_57);
            control_274_57 <= (control_274_56);
            control_274_56 <= (control_274_55);
            control_274_55 <= (control_274_54);
            control_274_54 <= (control_274_53);
            control_274_53 <= (control_274_52);
            control_274_52 <= (control_274_51);
            control_274_51 <= (control_274_50);
            control_274_50 <= (control_274_49);
            control_274_49 <= (control_274_48);
            control_274_48 <= (control_274_47);
            control_274_47 <= (control_274_46);
            control_274_46 <= (control_274_45);
            control_274_45 <= (control_274_44);
            control_274_44 <= (control_274_43);
            control_274_43 <= (control_274_42);
            control_274_42 <= (control_274_41);
            control_274_41 <= (control_274_40);
            control_274_40 <= (control_274_39);
            control_274_39 <= (control_274_38);
            control_274_38 <= (control_274_37);
            control_274_37 <= (control_274_36);
            control_274_36 <= (control_274_35);
            control_274_35 <= (control_274_34);
            control_274_34 <= (control_274_33);
            control_274_33 <= (control_274_32);
            control_274_32 <= (control_274_31);
            control_274_31 <= (control_274_30);
            control_274_30 <= (control_274_29);
            control_274_29 <= (control_274_28);
            control_274_28 <= (control_274_27);
            control_274_27 <= (control_274_26);
            control_274_26 <= (control_274_25);
            control_274_25 <= (control_274_24);
            control_274_24 <= (control_274_23);
            control_274_23 <= (control_274_22);
            control_274_22 <= (control_274_21);
            control_274_21 <= (control_274_20);
            control_274_20 <= (control_274_19);
            control_274_19 <= (control_274_18);
            control_274_18 <= (control_274_17);
            control_274_17 <= (control_274_16);
            control_274_16 <= (control_274_15);
            control_274_15 <= (control_274_14);
            control_274_14 <= (control_274_13);
            control_274_13 <= (control_274_12);
            control_274_12 <= (control_274_11);
            control_274_11 <= (control_274_10);
            control_274_10 <= (control_274_9);
            control_274_9 <= (control_274_8);
            control_274_8 <= (control_274_7);
            control_274_7 <= (control_274_6);
            control_274_6 <= (control_274_5);
            control_274_5 <= (control_274_4);
            control_274_4 <= (control_274_3);
            control_274_3 <= (control_274_2);
            control_274_2 <= (control_274_1);
            control_274_1 <= (control_274_start);
            input_key_274_follow <= (input_key_274);
            input_in_274_follow <= (input_in_274);
            lookup_sbox_0_output <= ((lookup_sbox_0_enable)?(sbox_0[(lookup_sbox_0_0)]):(lookup_sbox_0_output));
            lookup_sbox_1_output <= ((lookup_sbox_1_enable)?(sbox_1[(lookup_sbox_1_0)]):(lookup_sbox_1_output));
            lookup_sbox_2_output <= ((lookup_sbox_2_enable)?(sbox_2[(lookup_sbox_2_0)]):(lookup_sbox_2_output));
            lookup_sbox_3_output <= ((lookup_sbox_3_enable)?(sbox_3[(lookup_sbox_3_0)]):(lookup_sbox_3_output));
            lookup_sbox_4_output <= ((lookup_sbox_4_enable)?(sbox_4[(lookup_sbox_4_0)]):(lookup_sbox_4_output));
            lookup_sbox_5_output <= ((lookup_sbox_5_enable)?(sbox_5[(lookup_sbox_5_0)]):(lookup_sbox_5_output));
            lookup_sbox_6_output <= ((lookup_sbox_6_enable)?(sbox_6[(lookup_sbox_6_0)]):(lookup_sbox_6_output));
            lookup_sbox_7_output <= ((lookup_sbox_7_enable)?(sbox_7[(lookup_sbox_7_0)]):(lookup_sbox_7_output));
            lookup_sbox_8_output <= ((lookup_sbox_8_enable)?(sbox_8[(lookup_sbox_8_0)]):(lookup_sbox_8_output));
            lookup_sbox_9_output <= ((lookup_sbox_9_enable)?(sbox_9[(lookup_sbox_9_0)]):(lookup_sbox_9_output));
            lookup_sbox_10_output <= ((lookup_sbox_10_enable)?(sbox_10[(lookup_sbox_10_0)]):(lookup_sbox_10_output));
            lookup_sbox_11_output <= ((lookup_sbox_11_enable)?(sbox_11[(lookup_sbox_11_0)]):(lookup_sbox_11_output));
            lookup_sbox_12_output <= ((lookup_sbox_12_enable)?(sbox_12[(lookup_sbox_12_0)]):(lookup_sbox_12_output));
            lookup_sbox_13_output <= ((lookup_sbox_13_enable)?(sbox_13[(lookup_sbox_13_0)]):(lookup_sbox_13_output));
            lookup_sbox_14_output <= ((lookup_sbox_14_enable)?(sbox_14[(lookup_sbox_14_0)]):(lookup_sbox_14_output));
            lookup_sbox_15_output <= ((lookup_sbox_15_enable)?(sbox_15[(lookup_sbox_15_0)]):(lookup_sbox_15_output));
            startfollow <= (start);
        end
endmodule // end of module AES128_encrypt
